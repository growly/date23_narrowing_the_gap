`define  n 32
`define max_size 30

module dual_port_ram(clk, we1, we2, addr1, addr2, data1, data2, out1, out2);
parameter ADDR_WIDTH = 12;
parameter DATA_WIDTH = 32;
input clk;
input we1, we2;
input [ADDR_WIDTH-1:0] addr1, addr2;
input [DATA_WIDTH-1:0] data1, data2;
output reg [DATA_WIDTH-1:0] out1, out2;
reg [DATA_WIDTH-1:0] RAM [(1<<ADDR_WIDTH)-1:0];
always @(posedge clk)
begin
    if (we1)
            RAM[addr1] <= data1;
    if (we2)
            RAM[addr2] <= data2;
    out1 <= RAM[addr1];
    out2 <= RAM[addr2];
end
endmodule


//
// Generated by Bluespec Compiler, version 2009.11.beta2 (build 18693, 2009-11-24)
//
// On Tue Jun  8 18:43:40 EDT 2010
//
//
// Ports:
// Name                         I/O  size props
// wciS0_SResp                    O     2 reg
// wciS0_SData                    O    32 reg
// wciS0_SThreadBusy              O     1
// wciS0_SFlag                    O     2
// wsiS1_SThreadBusy              O     1
// wsiS1_SReset_n                 O     1
// wsiM1_MCmd                     O     3
// wsiM1_MReqLast                 O     1
// wsiM1_MBurstPrecise            O     1
// wsiM1_MBurstLength             O    12
// wsiM1_MData                    O   256 reg
// wsiM1_MByteEn                  O    32 reg
// wsiM1_MReqInfo                 O     8
// wsiM1_MReset_n                 O     1
// wmemiM_MCmd                    O     3 reg
// wmemiM_MReqLast                O     1 reg
// wmemiM_MAddr                   O    36 reg
// wmemiM_MBurstLength            O    12 reg
// wmemiM_MDataValid              O     1 reg
// wmemiM_MDataLast               O     1 reg
// wmemiM_MData                   O   128 reg
// wmemiM_MDataByteEn             O    16 reg
// wmemiM_MReset_n                O     1
// wciS0_Clk                      I     1 clock
// wciS0_MReset_n                 I     1 reset
// wciS0_MCmd                     I     3
// wciS0_MAddrSpace               I     1
// wciS0_MByteEn                  I     4
// wciS0_MAddr                    I    20
// wciS0_MData                    I    32
// wciS0_MFlag                    I     2 unused
// wsiS1_MCmd                     I     3
// wsiS1_MBurstLength             I    12
// wsiS1_MData                    I   256
// wsiS1_MByteEn                  I    32
// wsiS1_MReqInfo                 I     8
// wmemiM_SResp                   I     2
// wmemiM_SData                   I   128
// wsiS1_MReqLast                 I     1
// wsiS1_MBurstPrecise            I     1
// wsiS1_MReset_n                 I     1 reg
// wsiM1_SThreadBusy              I     1 reg
// wsiM1_SReset_n                 I     1 reg
// wmemiM_SRespLast               I     1
// wmemiM_SCmdAccept              I     1
// wmemiM_SDataAccept             I     1
//
// No combinational paths from inputs to outputs
//
//



module mkDelayWorker32B(wciS0_Clk,
			wciS0_MReset_n,

			wciS0_MCmd,

			wciS0_MAddrSpace,

			wciS0_MByteEn,

			wciS0_MAddr,

			wciS0_MData,

			wciS0_SResp,

			wciS0_SData,

			wciS0_SThreadBusy,

			wciS0_SFlag,

			wciS0_MFlag,

			wsiS1_MCmd,

			wsiS1_MReqLast,

			wsiS1_MBurstPrecise,

			wsiS1_MBurstLength,

			wsiS1_MData,

			wsiS1_MByteEn,

			wsiS1_MReqInfo,

			wsiS1_SThreadBusy,

			wsiS1_SReset_n,

			wsiS1_MReset_n,

			wsiM1_MCmd,

			wsiM1_MReqLast,

			wsiM1_MBurstPrecise,

			wsiM1_MBurstLength,

			wsiM1_MData,

			wsiM1_MByteEn,

			wsiM1_MReqInfo,

			wsiM1_SThreadBusy,

			wsiM1_MReset_n,

			wsiM1_SReset_n,

			wmemiM_MCmd,

			wmemiM_MReqLast,

			wmemiM_MAddr,

			wmemiM_MBurstLength,

			wmemiM_MDataValid,

			wmemiM_MDataLast,

			wmemiM_MData,

			wmemiM_MDataByteEn,

			wmemiM_SResp,

			wmemiM_SRespLast,

			wmemiM_SData,

			wmemiM_SCmdAccept,

			wmemiM_SDataAccept,

			wmemiM_MReset_n,
			
			prevent_hanging_nodes);
  parameter [31 : 0] dlyCtrlInit = 32'b00000000000000000000000000000000;
  input  wciS0_Clk;
  input  wciS0_MReset_n;

  // action method wciS0_mCmd
  input  [2 : 0] wciS0_MCmd;

  // action method wciS0_mAddrSpace
  input  wciS0_MAddrSpace;

  // action method wciS0_mByteEn
  input  [3 : 0] wciS0_MByteEn;

  // action method wciS0_mAddr
  input  [19 : 0] wciS0_MAddr;

  // action method wciS0_mData
  input  [31 : 0] wciS0_MData;

  // value method wciS0_sResp
  output [1 : 0] wciS0_SResp;

  // value method wciS0_sData
  output [31 : 0] wciS0_SData;

  // value method wciS0_sThreadBusy
  output wciS0_SThreadBusy;

  // value method wciS0_sFlag
  output [1 : 0] wciS0_SFlag;

  // action method wciS0_mFlag
  input  [1 : 0] wciS0_MFlag;

  // action method wsiS1_mCmd
  input  [2 : 0] wsiS1_MCmd;

  // action method wsiS1_mReqLast
  input  wsiS1_MReqLast;

  // action method wsiS1_mBurstPrecise
  input  wsiS1_MBurstPrecise;

  // action method wsiS1_mBurstLength
  input  [11 : 0] wsiS1_MBurstLength;

  // action method wsiS1_mData
  input  [255 : 0] wsiS1_MData;

  // action method wsiS1_mByteEn
  input  [31 : 0] wsiS1_MByteEn;

  // action method wsiS1_mReqInfo
  input  [7 : 0] wsiS1_MReqInfo;

  // action method wsiS1_mDataInfo

  // value method wsiS1_sThreadBusy
  output wsiS1_SThreadBusy;

  // value method wsiS1_sReset_n
  output wsiS1_SReset_n;

  // action method wsiS1_mReset_n
  input  wsiS1_MReset_n;

  // value method wsiM1_mCmd
  output [2 : 0] wsiM1_MCmd;

  // value method wsiM1_mReqLast
  output wsiM1_MReqLast;

  // value method wsiM1_mBurstPrecise
  output wsiM1_MBurstPrecise;

  // value method wsiM1_mBurstLength
  output [11 : 0] wsiM1_MBurstLength;

  // value method wsiM1_mData
  output [255 : 0] wsiM1_MData;

  // value method wsiM1_mByteEn
  output [31 : 0] wsiM1_MByteEn;

  // value method wsiM1_mReqInfo
  output [7 : 0] wsiM1_MReqInfo;

  // value method wsiM1_mDataInfo

  // action method wsiM1_sThreadBusy
  input  wsiM1_SThreadBusy;

  // value method wsiM1_mReset_n
  output wsiM1_MReset_n;

  // action method wsiM1_sReset_n
  input  wsiM1_SReset_n;

  // value method wmemiM_mCmd
  output [2 : 0] wmemiM_MCmd;

  // value method wmemiM_mReqLast
  output wmemiM_MReqLast;

  // value method wmemiM_mAddr
  output [35 : 0] wmemiM_MAddr;

  // value method wmemiM_mBurstLength
  output [11 : 0] wmemiM_MBurstLength;

  // value method wmemiM_mDataValid
  output wmemiM_MDataValid;

  // value method wmemiM_mDataLast
  output wmemiM_MDataLast;

  // value method wmemiM_mData
  output [127 : 0] wmemiM_MData;

  // value method wmemiM_mDataByteEn
  output [15 : 0] wmemiM_MDataByteEn;

  // action method wmemiM_sResp
  input  [1 : 0] wmemiM_SResp;

  // action method wmemiM_sRespLast
  input  wmemiM_SRespLast;

  // action method wmemiM_sData
  input  [127 : 0] wmemiM_SData;

  // action method wmemiM_sCmdAccept
  input  wmemiM_SCmdAccept;

  // action method wmemiM_sDataAccept
  input  wmemiM_SDataAccept;

  // value method wmemiM_mReset_n
  output wmemiM_MReset_n;
  
  output prevent_hanging_nodes;

  // Hanging node logic
  
  
  
  wire dummy1;
  wire dummy2;
  wire dummy3;
  wire dummy4;
  wire dummy5;
  wire dummy6;
  wire dummy7;
  wire dummy8;
  wire dummy9;
  assign dummy1 = &mesgRF_memory__DOB;
  assign dummy2 = &mesgWF_memory__DOB;
  assign dummy3 = &metaRF__D_OUT;
  assign dummy4 = &metaWF__D_OUT ;
  assign dummy5 = &wci_reqF__D_OUT;
  assign dummy6 = &wide16Fa__D_OUT;
  assign dummy7 = &wide16Fb__D_OUT;
  assign dummy8 = &wmemi_respF__D_OUT;
  assign dummy9 = &wsiS_reqFifo__D_OUT;
  
  wire prevent_hang_wire;
  assign prevent_hang_wire =  dummy1 & dummy2 & dummy3 & dummy4 &dummy5 & dummy6 & dummy7 & dummy8 & dummy9;
  assign prevent_hanging_nodes = prevent_hang_wire;

  // signals for module outputs
  wire [255 : 0] wsiM1_MData;
  wire [127 : 0] wmemiM_MData;
  wire [35 : 0] wmemiM_MAddr;
  wire [31 : 0] wciS0_SData, wsiM1_MByteEn;
  wire [15 : 0] wmemiM_MDataByteEn;
  wire [11 : 0] wmemiM_MBurstLength, wsiM1_MBurstLength;
  wire [7 : 0] wsiM1_MReqInfo;
  wire [2 : 0] wmemiM_MCmd, wsiM1_MCmd;
  wire [1 : 0] wciS0_SFlag, wciS0_SResp;
  wire wciS0_SThreadBusy,
       wmemiM_MDataLast,
       wmemiM_MDataValid,
       wmemiM_MReqLast,
       wmemiM_MReset_n,
       wsiM1_MBurstPrecise,
       wsiM1_MReqLast,
       wsiM1_MReset_n,
       wsiS1_SReset_n,
       wsiS1_SThreadBusy;

  // inlined wires
  wire [312 : 0] wsiM_reqFifo_x_wire__wget, wsiS_wsiReq__wget;
  wire [255 : 0] mesgRF_wDataIn__wget,
		 mesgRF_wDataOut__wget,
		 mesgWF_wDataIn__wget,
		 mesgWF_wDataOut__wget,
		 wsi_Es_mData_w__wget;
  wire [145 : 0] wmemi_dhF_x_wire__wget;
  wire [130 : 0] wmemi_wmemiResponse__wget;
  wire [127 : 0] wmemi_Em_sData_w__wget;
  wire [95 : 0] wsiM_extStatusW__wget, wsiS_extStatusW__wget;
  wire [59 : 0] wci_wciReq__wget;
  wire [51 : 0] wmemi_reqF_x_wire__wget;
  wire [33 : 0] wci_respF_x_wire__wget;
  wire [31 : 0] wci_Es_mData_w__wget, wsi_Es_mByteEn_w__wget;
  wire [19 : 0] dlyWordsStored_acc_v1__wget,
		dlyWordsStored_acc_v2__wget,
		wci_Es_mAddr_w__wget;
  wire [11 : 0] wsi_Es_mBurstLength_w__wget;
  wire [7 : 0] dlyReadCredit_acc_v1__wget,
	       dlyReadCredit_acc_v2__wget,
	       wsi_Es_mReqInfo_w__wget;
  wire [3 : 0] wci_Es_mByteEn_w__wget;
  wire [2 : 0] wci_Es_mCmd_w__wget, wci_wEdge__wget, wsi_Es_mCmd_w__wget;
  wire [1 : 0] wmemi_Em_sResp_w__wget;
  wire dlyReadCredit_acc_v1__whas,
       dlyReadCredit_acc_v2__whas,
       dlyWordsStored_acc_v1__whas,
       dlyWordsStored_acc_v2__whas,
       mesgRF_pwDequeue__whas,
       mesgRF_pwEnqueue__whas,
       mesgRF_wDataIn__whas,
       mesgRF_wDataOut__whas,
       mesgWF_pwDequeue__whas,
       mesgWF_pwEnqueue__whas,
       mesgWF_wDataIn__whas,
       mesgWF_wDataOut__whas,
       wci_Es_mAddrSpace_w__wget,
       wci_Es_mAddrSpace_w__whas,
       wci_Es_mAddr_w__whas,
       wci_Es_mByteEn_w__whas,
       wci_Es_mCmd_w__whas,
       wci_Es_mData_w__whas,
       wci_ctlAckReg_1__wget,
       wci_ctlAckReg_1__whas,
       wci_reqF_r_clr__whas,
       wci_reqF_r_deq__whas,
       wci_reqF_r_enq__whas,
       wci_respF_dequeueing__whas,
       wci_respF_enqueueing__whas,
       wci_respF_x_wire__whas,
       wci_sFlagReg_1__wget,
       wci_sFlagReg_1__whas,
       wci_sThreadBusy_pw__whas,
       wci_wEdge__whas,
       wci_wciReq__whas,
       wci_wci_cfrd_pw__whas,
       wci_wci_cfwr_pw__whas,
       wci_wci_ctrl_pw__whas,
       wmemi_Em_sData_w__whas,
       wmemi_Em_sRespLast_w__whas,
       wmemi_Em_sResp_w__whas,
       wmemi_dhF_dequeueing__whas,
       wmemi_dhF_enqueueing__whas,
       wmemi_dhF_x_wire__whas,
       wmemi_operateD_1__wget,
       wmemi_operateD_1__whas,
       wmemi_peerIsReady_1__wget,
       wmemi_peerIsReady_1__whas,
       wmemi_reqF_dequeueing__whas,
       wmemi_reqF_enqueueing__whas,
       wmemi_reqF_x_wire__whas,
       wmemi_sCmdAccept_w__wget,
       wmemi_sCmdAccept_w__whas,
       wmemi_sDataAccept_w__wget,
       wmemi_sDataAccept_w__whas,
       wmemi_wmemiResponse__whas,
       wsiM_operateD_1__wget,
       wsiM_operateD_1__whas,
       wsiM_peerIsReady_1__wget,
       wsiM_peerIsReady_1__whas,
       wsiM_reqFifo_dequeueing__whas,
       wsiM_reqFifo_enqueueing__whas,
       wsiM_reqFifo_x_wire__whas,
       wsiM_sThreadBusy_pw__whas,
       wsiS_operateD_1__wget,
       wsiS_operateD_1__whas,
       wsiS_peerIsReady_1__wget,
       wsiS_peerIsReady_1__whas,
       wsiS_reqFifo_r_clr__whas,
       wsiS_reqFifo_r_deq__whas,
       wsiS_reqFifo_r_enq__whas,
       wsiS_wsiReq__whas,
       wsi_Es_mBurstLength_w__whas,
       wsi_Es_mBurstPrecise_w__whas,
       wsi_Es_mByteEn_w__whas,
       wsi_Es_mCmd_w__whas,
       wsi_Es_mDataInfo_w__whas,
       wsi_Es_mData_w__whas,
       wsi_Es_mReqInfo_w__whas,
       wsi_Es_mReqLast_w__whas;

  // register abortCount
  reg [31 : 0] abortCount;
  wire [31 : 0] abortCount__D_IN;
  wire abortCount__EN;

  // register blockDelayWrite
  reg blockDelayWrite;
  wire blockDelayWrite__D_IN, blockDelayWrite__EN;

  // register bytesRead
  reg [31 : 0] bytesRead;
  wire [31 : 0] bytesRead__D_IN;
  wire bytesRead__EN;

  // register bytesWritten
  reg [31 : 0] bytesWritten;
  wire [31 : 0] bytesWritten__D_IN;
  wire bytesWritten__EN;

  // register cyclesPassed
  reg [31 : 0] cyclesPassed;
  wire [31 : 0] cyclesPassed__D_IN;
  wire cyclesPassed__EN;

  // register dlyCtrl
  reg [31 : 0] dlyCtrl;
  wire [31 : 0] dlyCtrl__D_IN;
  wire dlyCtrl__EN;

  // register dlyHoldoffBytes
  reg [31 : 0] dlyHoldoffBytes;
  wire [31 : 0] dlyHoldoffBytes__D_IN;
  wire dlyHoldoffBytes__EN;

  // register dlyHoldoffCycles
  reg [31 : 0] dlyHoldoffCycles;
  wire [31 : 0] dlyHoldoffCycles__D_IN;
  wire dlyHoldoffCycles__EN;

  // register dlyRAG
  reg [19 : 0] dlyRAG;
  wire [19 : 0] dlyRAG__D_IN;
  wire dlyRAG__EN;

  // register dlyReadCredit_value
  reg [7 : 0] dlyReadCredit_value;
  wire [7 : 0] dlyReadCredit_value__D_IN;
  wire dlyReadCredit_value__EN;

  // register dlyWAG
  reg [19 : 0] dlyWAG;
  wire [19 : 0] dlyWAG__D_IN;
  wire dlyWAG__EN;

  // register dlyWordsStored_value
  reg [19 : 0] dlyWordsStored_value;
  wire [19 : 0] dlyWordsStored_value__D_IN;
  wire dlyWordsStored_value__EN;

  // register doAbort
  reg doAbort;
  wire doAbort__D_IN, doAbort__EN;

  // register endOfMessage
  reg endOfMessage;
  wire endOfMessage__D_IN, endOfMessage__EN;

  // register errCount // jluu removed because never used
//  reg [255 : 0] errCount;
//  wire [255 : 0] errCount__D_IN;
//  wire errCount__EN;

  // register impreciseBurst
  reg impreciseBurst;
  reg impreciseBurst__D_IN;
  wire impreciseBurst__EN;

  // register mesgLength
  reg [14 : 0] mesgLength;
  reg [14 : 0] mesgLength__D_IN;
  wire mesgLength__EN;

  // register mesgLengthSoFar
  reg [13 : 0] mesgLengthSoFar;
  wire [13 : 0] mesgLengthSoFar__D_IN;
  wire mesgLengthSoFar__EN;

  // register mesgRF_rCache
  reg [267 : 0] mesgRF_rCache;
  wire [267 : 0] mesgRF_rCache__D_IN;
  wire mesgRF_rCache__EN;

  // register mesgRF_rRdPtr
  reg [10 : 0] mesgRF_rRdPtr;
  wire [10 : 0] mesgRF_rRdPtr__D_IN;
  wire mesgRF_rRdPtr__EN;

  // register mesgRF_rWrPtr
  reg [10 : 0] mesgRF_rWrPtr;
  wire [10 : 0] mesgRF_rWrPtr__D_IN;
  wire mesgRF_rWrPtr__EN;

  // register mesgRdCount
  reg [31 : 0] mesgRdCount;
  wire [31 : 0] mesgRdCount__D_IN;
  wire mesgRdCount__EN;

  // register mesgReqValid
  reg mesgReqValid;
  wire mesgReqValid__D_IN, mesgReqValid__EN;

  // register mesgWF_rCache
  reg [267 : 0] mesgWF_rCache;
  wire [267 : 0] mesgWF_rCache__D_IN;
  wire mesgWF_rCache__EN;

  // register mesgWF_rRdPtr
  reg [10 : 0] mesgWF_rRdPtr;
  wire [10 : 0] mesgWF_rRdPtr__D_IN;
  wire mesgWF_rRdPtr__EN;

  // register mesgWF_rWrPtr
  reg [10 : 0] mesgWF_rWrPtr;
  wire [10 : 0] mesgWF_rWrPtr__D_IN;
  wire mesgWF_rWrPtr__EN;

  // register mesgWtCount
  reg [31 : 0] mesgWtCount;
  wire [31 : 0] mesgWtCount__D_IN;
  wire mesgWtCount__EN;

  // register opcode
  reg [8 : 0] opcode;
  reg [8 : 0] opcode__D_IN;
  wire opcode__EN;

  // register preciseBurst
  reg preciseBurst;
  reg preciseBurst__D_IN;
  wire preciseBurst__EN;

  // register rdSerAddr
  reg [31 : 0] rdSerAddr;
  wire [31 : 0] rdSerAddr__D_IN;
  wire rdSerAddr__EN;

  // register rdSerEmpty
  reg rdSerEmpty;
  wire rdSerEmpty__D_IN, rdSerEmpty__EN;

  // register rdSerMeta
  reg [31 : 0] rdSerMeta;
  wire [31 : 0] rdSerMeta__D_IN;
  wire rdSerMeta__EN;

  // register rdSerPos
  reg [1 : 0] rdSerPos;
  wire [1 : 0] rdSerPos__D_IN;
  wire rdSerPos__EN;

  // register rdSerStage
  reg [31 : 0] rdSerStage;
  wire [31 : 0] rdSerStage__D_IN;
  wire rdSerStage__EN;

  // register rdSerStage_1
  reg [31 : 0] rdSerStage_1;
  wire [31 : 0] rdSerStage_1__D_IN;
  wire rdSerStage_1__EN;

  // register rdSerStage_2
  reg [31 : 0] rdSerStage_2;
  wire [31 : 0] rdSerStage_2__D_IN;
  wire rdSerStage_2__EN;

  // register rdSerStage_3
  reg [31 : 0] rdSerStage_3;
  wire [31 : 0] rdSerStage_3__D_IN;
  wire rdSerStage_3__EN;

  // register rdSerUnroll
  reg [15 : 0] rdSerUnroll;
  wire [15 : 0] rdSerUnroll__D_IN;
  wire rdSerUnroll__EN;

  // register rdSyncWord
  reg rdSyncWord;
  reg rdSyncWord__D_IN;
  wire rdSyncWord__EN;

  // register readMeta
  reg [31 : 0] readMeta;
  wire [31 : 0] readMeta__D_IN;
  wire readMeta__EN;

  // register readyToPush
  reg readyToPush;
  reg readyToPush__D_IN;
  wire readyToPush__EN;

  // register readyToRequest
  reg readyToRequest;
  wire readyToRequest__D_IN, readyToRequest__EN;

  // register unrollCnt
  reg [15 : 0] unrollCnt;
  wire [15 : 0] unrollCnt__D_IN;
  wire unrollCnt__EN;

  // register valExpect
//  reg [255 : 0] valExpect;
//  wire [255 : 0] valExpect__D_IN;
//  wire valExpect__EN;

  // register wci_cEdge
  reg [2 : 0] wci_cEdge;
  wire [2 : 0] wci_cEdge__D_IN;
  wire wci_cEdge__EN;

  // register wci_cState
  reg [2 : 0] wci_cState;
  wire [2 : 0] wci_cState__D_IN;
  wire wci_cState__EN;

  // register wci_ctlAckReg
  reg wci_ctlAckReg;
  wire wci_ctlAckReg__D_IN, wci_ctlAckReg__EN;

  // register wci_ctlOpActive
  reg wci_ctlOpActive;
  wire wci_ctlOpActive__D_IN, wci_ctlOpActive__EN;

  // register wci_illegalEdge
  reg wci_illegalEdge;
  wire wci_illegalEdge__D_IN, wci_illegalEdge__EN;

  // register wci_nState
  reg [2 : 0] wci_nState;
  reg [2 : 0] wci_nState__D_IN;
  wire wci_nState__EN;

  // register wci_reqF_countReg
  reg [1 : 0] wci_reqF_countReg;
  wire [1 : 0] wci_reqF_countReg__D_IN;
  wire wci_reqF_countReg__EN;

  // register wci_respF_c_r
  reg [1 : 0] wci_respF_c_r;
  wire [1 : 0] wci_respF_c_r__D_IN;
  wire wci_respF_c_r__EN;

  // register wci_respF_q_0
  reg [33 : 0] wci_respF_q_0;
  reg [33 : 0] wci_respF_q_0__D_IN;
  wire wci_respF_q_0__EN;

  // register wci_respF_q_1
  reg [33 : 0] wci_respF_q_1;
  reg [33 : 0] wci_respF_q_1__D_IN;
  wire wci_respF_q_1__EN;

  // register wci_sFlagReg
  reg wci_sFlagReg;
  wire wci_sFlagReg__D_IN, wci_sFlagReg__EN;

  // register wci_sThreadBusy_d
  reg wci_sThreadBusy_d;
  wire wci_sThreadBusy_d__D_IN, wci_sThreadBusy_d__EN;

  // register wmemiRdReq
  reg [31 : 0] wmemiRdReq;
  wire [31 : 0] wmemiRdReq__D_IN;
  wire wmemiRdReq__EN;

  // register wmemiRdResp
  reg [31 : 0] wmemiRdResp;
  wire [31 : 0] wmemiRdResp__D_IN;
  wire wmemiRdResp__EN;

  // register wmemiWrReq
  reg [31 : 0] wmemiWrReq;
  wire [31 : 0] wmemiWrReq__D_IN;
  wire wmemiWrReq__EN;

  // register wmemi_busyWithMessage
  reg wmemi_busyWithMessage;
  wire wmemi_busyWithMessage__D_IN, wmemi_busyWithMessage__EN;

  // register wmemi_dhF_c_r
  reg [1 : 0] wmemi_dhF_c_r;
  wire [1 : 0] wmemi_dhF_c_r__D_IN;
  wire wmemi_dhF_c_r__EN;

  // register wmemi_dhF_q_0
  reg [145 : 0] wmemi_dhF_q_0;
  reg [145 : 0] wmemi_dhF_q_0__D_IN;
  wire wmemi_dhF_q_0__EN;

  // register wmemi_dhF_q_1
  reg [145 : 0] wmemi_dhF_q_1;
  reg [145 : 0] wmemi_dhF_q_1__D_IN;
  wire wmemi_dhF_q_1__EN;

  // register wmemi_errorSticky
  reg wmemi_errorSticky;
  wire wmemi_errorSticky__D_IN, wmemi_errorSticky__EN;

  // register wmemi_operateD
  reg wmemi_operateD;
  wire wmemi_operateD__D_IN, wmemi_operateD__EN;

  // register wmemi_peerIsReady
  reg wmemi_peerIsReady;
  wire wmemi_peerIsReady__D_IN, wmemi_peerIsReady__EN;

  // register wmemi_reqF_c_r
  reg [1 : 0] wmemi_reqF_c_r;
  wire [1 : 0] wmemi_reqF_c_r__D_IN;
  wire wmemi_reqF_c_r__EN;

  // register wmemi_reqF_q_0
  reg [51 : 0] wmemi_reqF_q_0;
  reg [51 : 0] wmemi_reqF_q_0__D_IN;
  wire wmemi_reqF_q_0__EN;

  // register wmemi_reqF_q_1
  reg [51 : 0] wmemi_reqF_q_1;
  reg [51 : 0] wmemi_reqF_q_1__D_IN;
  wire wmemi_reqF_q_1__EN;

  // register wmemi_statusR
  reg [7 : 0] wmemi_statusR;
  wire [7 : 0] wmemi_statusR__D_IN;
  wire wmemi_statusR__EN;

  // register wmemi_trafficSticky
  reg wmemi_trafficSticky;
  wire wmemi_trafficSticky__D_IN, wmemi_trafficSticky__EN;

  // register wrtDutyCount
  reg [2 : 0] wrtDutyCount;
  wire [2 : 0] wrtDutyCount__D_IN;
  wire wrtDutyCount__EN;

  // register wrtSerAddr
  reg [31 : 0] wrtSerAddr;
  wire [31 : 0] wrtSerAddr__D_IN;
  wire wrtSerAddr__EN;

  // register wrtSerMeta
  reg [31 : 0] wrtSerMeta;
  wire [31 : 0] wrtSerMeta__D_IN;
  wire wrtSerMeta__EN;

  // register wrtSerPos
  reg [1 : 0] wrtSerPos;
  wire [1 : 0] wrtSerPos__D_IN;
  wire wrtSerPos__EN;

  // register wrtSerStage
  reg [31 : 0] wrtSerStage;
  wire [31 : 0] wrtSerStage__D_IN;
  wire wrtSerStage__EN;

  // register wrtSerStage_1
  reg [31 : 0] wrtSerStage_1;
  wire [31 : 0] wrtSerStage_1__D_IN;
  wire wrtSerStage_1__EN;

  // register wrtSerStage_2
  reg [31 : 0] wrtSerStage_2;
  wire [31 : 0] wrtSerStage_2__D_IN;
  wire wrtSerStage_2__EN;

  // register wrtSerStage_3
  reg [31 : 0] wrtSerStage_3;
  wire [31 : 0] wrtSerStage_3__D_IN;
  wire wrtSerStage_3__EN;

  // register wrtSerUnroll
  reg [15 : 0] wrtSerUnroll;
  wire [15 : 0] wrtSerUnroll__D_IN;
  wire wrtSerUnroll__EN;

  // register wsiM_burstKind
  reg [1 : 0] wsiM_burstKind;
  wire [1 : 0] wsiM_burstKind__D_IN;
  wire wsiM_burstKind__EN;

  // register wsiM_errorSticky
  reg wsiM_errorSticky;
  wire wsiM_errorSticky__D_IN, wsiM_errorSticky__EN;

  // register wsiM_iMesgCount
  reg [31 : 0] wsiM_iMesgCount;
  wire [31 : 0] wsiM_iMesgCount__D_IN;
  wire wsiM_iMesgCount__EN;

  // register wsiM_operateD
  reg wsiM_operateD;
  wire wsiM_operateD__D_IN, wsiM_operateD__EN;

  // register wsiM_pMesgCount
  reg [31 : 0] wsiM_pMesgCount;
  wire [31 : 0] wsiM_pMesgCount__D_IN;
  wire wsiM_pMesgCount__EN;

  // register wsiM_peerIsReady
  reg wsiM_peerIsReady;
  wire wsiM_peerIsReady__D_IN, wsiM_peerIsReady__EN;

  // register wsiM_reqFifo_c_r
  reg [1 : 0] wsiM_reqFifo_c_r;
  wire [1 : 0] wsiM_reqFifo_c_r__D_IN;
  wire wsiM_reqFifo_c_r__EN;

  // register wsiM_reqFifo_q_0
  reg [312 : 0] wsiM_reqFifo_q_0;
  reg [312 : 0] wsiM_reqFifo_q_0__D_IN;
  wire wsiM_reqFifo_q_0__EN;

  // register wsiM_reqFifo_q_1
  reg [312 : 0] wsiM_reqFifo_q_1;
  reg [312 : 0] wsiM_reqFifo_q_1__D_IN;
  wire wsiM_reqFifo_q_1__EN;

  // register wsiM_sThreadBusy_d
  reg wsiM_sThreadBusy_d;
  wire wsiM_sThreadBusy_d__D_IN, wsiM_sThreadBusy_d__EN;

  // register wsiM_statusR
  reg [7 : 0] wsiM_statusR;
  wire [7 : 0] wsiM_statusR__D_IN;
  wire wsiM_statusR__EN;

  // register wsiM_tBusyCount
  reg [31 : 0] wsiM_tBusyCount;
  wire [31 : 0] wsiM_tBusyCount__D_IN;
  wire wsiM_tBusyCount__EN;

  // register wsiM_trafficSticky
  reg wsiM_trafficSticky;
  wire wsiM_trafficSticky__D_IN, wsiM_trafficSticky__EN;

  // register wsiS_burstKind
  reg [1 : 0] wsiS_burstKind;
  wire [1 : 0] wsiS_burstKind__D_IN;
  wire wsiS_burstKind__EN;

  // register wsiS_errorSticky
  reg wsiS_errorSticky;
  wire wsiS_errorSticky__D_IN, wsiS_errorSticky__EN;

  // register wsiS_iMesgCount
  reg [31 : 0] wsiS_iMesgCount;
  wire [31 : 0] wsiS_iMesgCount__D_IN;
  wire wsiS_iMesgCount__EN;

  // register wsiS_operateD
  reg wsiS_operateD;
  wire wsiS_operateD__D_IN, wsiS_operateD__EN;

  // register wsiS_pMesgCount
  reg [31 : 0] wsiS_pMesgCount;
  wire [31 : 0] wsiS_pMesgCount__D_IN;
  wire wsiS_pMesgCount__EN;

  // register wsiS_peerIsReady
  reg wsiS_peerIsReady;
  wire wsiS_peerIsReady__D_IN, wsiS_peerIsReady__EN;

  // register wsiS_reqFifo_countReg
  reg [1 : 0] wsiS_reqFifo_countReg;
  wire [1 : 0] wsiS_reqFifo_countReg__D_IN;
  wire wsiS_reqFifo_countReg__EN;

  // register wsiS_statusR
  reg [7 : 0] wsiS_statusR;
  wire [7 : 0] wsiS_statusR__D_IN;
  wire wsiS_statusR__EN;

  // register wsiS_tBusyCount
  reg [31 : 0] wsiS_tBusyCount;
  wire [31 : 0] wsiS_tBusyCount__D_IN;
  wire wsiS_tBusyCount__EN;

  // register wsiS_trafficSticky
  reg wsiS_trafficSticky;
  wire wsiS_trafficSticky__D_IN, wsiS_trafficSticky__EN;

  // register wsiWordsRemain
  reg [11 : 0] wsiWordsRemain;
  wire [11 : 0] wsiWordsRemain__D_IN;
  wire wsiWordsRemain__EN;

  // register zeroLengthMesg
  reg zeroLengthMesg;
  wire zeroLengthMesg__D_IN, zeroLengthMesg__EN;

  // ports of submodule mesgRF_memory
  wire [255 : 0] mesgRF_memory__DIA, mesgRF_memory__DIB, mesgRF_memory__DOB;
  wire [9 : 0] mesgRF_memory__ADDRA, mesgRF_memory__ADDRB;
  wire mesgRF_memory__ENA,
       mesgRF_memory__ENB,
       mesgRF_memory__WEA,
       mesgRF_memory__WEB;

  // ports of submodule mesgWF_memory
  wire [255 : 0] mesgWF_memory__DIA, mesgWF_memory__DIB, mesgWF_memory__DOB;
  wire [9 : 0] mesgWF_memory__ADDRA, mesgWF_memory__ADDRB;
  wire mesgWF_memory__ENA,
       mesgWF_memory__ENB,
       mesgWF_memory__WEA,
       mesgWF_memory__WEB;

  // ports of submodule metaRF
  reg [31 : 0] metaRF__D_IN;
  wire [31 : 0] metaRF__D_OUT;
  wire metaRF__CLR, metaRF__DEQ, metaRF__EMPTY_N, metaRF__ENQ, metaRF__FULL_N;

  // ports of submodule metaWF
  wire [31 : 0] metaWF__D_IN, metaWF__D_OUT;
  wire metaWF__CLR, metaWF__DEQ, metaWF__EMPTY_N, metaWF__ENQ, metaWF__FULL_N;

  // ports of submodule wci_isReset
  wire wci_isReset__VAL;

  // ports of submodule wci_reqF
  wire [59 : 0] wci_reqF__D_IN, wci_reqF__D_OUT;
  wire wci_reqF__CLR, wci_reqF__DEQ, wci_reqF__EMPTY_N, wci_reqF__ENQ;

  // ports of submodule wide16Fa
  wire [127 : 0] wide16Fa__D_IN, wide16Fa__D_OUT;
  wire wide16Fa__CLR,
       wide16Fa__DEQ,
       wide16Fa__EMPTY_N,
       wide16Fa__ENQ,
       wide16Fa__FULL_N;

  // ports of submodule wide16Fb
  wire [127 : 0] wide16Fb__D_IN, wide16Fb__D_OUT;
  wire wide16Fb__CLR,
       wide16Fb__DEQ,
       wide16Fb__EMPTY_N,
       wide16Fb__ENQ,
       wide16Fb__FULL_N;

  // ports of submodule wmemi_isReset
  wire wmemi_isReset__VAL;

  // ports of submodule wmemi_respF
  wire [130 : 0] wmemi_respF__D_IN, wmemi_respF__D_OUT;
  wire wmemi_respF__CLR,
       wmemi_respF__DEQ,
       wmemi_respF__EMPTY_N,
       wmemi_respF__ENQ,
       wmemi_respF__FULL_N;

  // ports of submodule wsiM_isReset
  wire wsiM_isReset__VAL;

  // ports of submodule wsiS_isReset
  wire wsiS_isReset__VAL;

  // ports of submodule wsiS_reqFifo
  wire [312 : 0] wsiS_reqFifo__D_IN, wsiS_reqFifo__D_OUT;
  wire wsiS_reqFifo__CLR,
       wsiS_reqFifo__DEQ,
       wsiS_reqFifo__EMPTY_N,
       wsiS_reqFifo__ENQ,
       wsiS_reqFifo__FULL_N;

  // rule scheduling signals
  wire CAN_FIRE_RL_cycles_passed_count,
       CAN_FIRE_RL_delay_read_req,
       CAN_FIRE_RL_delay_read_resp,
       CAN_FIRE_RL_delay_write_req,
       CAN_FIRE_RL_delay_write_unblock,
       CAN_FIRE_RL_dlyReadCredit_accumulate,
       CAN_FIRE_RL_dlyWordsStored_accumulate,
       CAN_FIRE_RL_mesgRF_portA,
       CAN_FIRE_RL_mesgRF_portB,
       CAN_FIRE_RL_mesgRF_portB_read_data,
       CAN_FIRE_RL_mesgWF_portA,
       CAN_FIRE_RL_mesgWF_portB,
       CAN_FIRE_RL_mesgWF_portB_read_data,
       CAN_FIRE_RL_operating_actions,
       CAN_FIRE_RL_rdSer_begin,
       CAN_FIRE_RL_rdSer_body,
       CAN_FIRE_RL_rdSer_sync,
       CAN_FIRE_RL_wci_Es_doAlways_Req,
       CAN_FIRE_RL_wci_cfrd,
       CAN_FIRE_RL_wci_cfwr,
       CAN_FIRE_RL_wci_ctlAckReg__dreg_update,
       CAN_FIRE_RL_wci_ctl_op_complete,
       CAN_FIRE_RL_wci_ctl_op_start,
       CAN_FIRE_RL_wci_ctrl_EiI,
       CAN_FIRE_RL_wci_ctrl_IsO,
       CAN_FIRE_RL_wci_ctrl_OrE,
       CAN_FIRE_RL_wci_reqF__updateLevelCounter,
       CAN_FIRE_RL_wci_reqF_enq,
       CAN_FIRE_RL_wci_request_decode,
       CAN_FIRE_RL_wci_respF_both,
       CAN_FIRE_RL_wci_respF_decCtr,
       CAN_FIRE_RL_wci_respF_deq,
       CAN_FIRE_RL_wci_respF_incCtr,
       CAN_FIRE_RL_wci_sFlagReg__dreg_update,
       CAN_FIRE_RL_wci_sThreadBusy_reg,
       CAN_FIRE_RL_wmemi_Em_doAlways,
       CAN_FIRE_RL_wmemi_dhF_both,
       CAN_FIRE_RL_wmemi_dhF_decCtr,
       CAN_FIRE_RL_wmemi_dhF_deq,
       CAN_FIRE_RL_wmemi_dhF_incCtr,
       CAN_FIRE_RL_wmemi_operateD__dreg_update,
       CAN_FIRE_RL_wmemi_peerIsReady__dreg_update,
       CAN_FIRE_RL_wmemi_reqF_both,
       CAN_FIRE_RL_wmemi_reqF_decCtr,
       CAN_FIRE_RL_wmemi_reqF_deq,
       CAN_FIRE_RL_wmemi_reqF_incCtr,
       CAN_FIRE_RL_wmemi_respAdvance,
       CAN_FIRE_RL_wmemi_update_statusR,
       CAN_FIRE_RL_wmrd_mesgBegin,
       CAN_FIRE_RL_wmrd_mesgBodyResponse,
       CAN_FIRE_RL_wmwt_doAbort,
       CAN_FIRE_RL_wmwt_mesgBegin,
       CAN_FIRE_RL_wmwt_messageFinalize,
       CAN_FIRE_RL_wmwt_messagePushImprecise,
       CAN_FIRE_RL_wmwt_messagePushPrecise,
       CAN_FIRE_RL_wmwt_requestPrecise,
       CAN_FIRE_RL_wrtSer_begin,
       CAN_FIRE_RL_wrtSer_body,
       CAN_FIRE_RL_wsiM_ext_status_assign,
       CAN_FIRE_RL_wsiM_inc_tBusyCount,
       CAN_FIRE_RL_wsiM_operateD__dreg_update,
       CAN_FIRE_RL_wsiM_peerIsReady__dreg_update,
       CAN_FIRE_RL_wsiM_reqFifo_both,
       CAN_FIRE_RL_wsiM_reqFifo_decCtr,
       CAN_FIRE_RL_wsiM_reqFifo_deq,
       CAN_FIRE_RL_wsiM_reqFifo_incCtr,
       CAN_FIRE_RL_wsiM_sThreadBusy_reg,
       CAN_FIRE_RL_wsiM_update_statusR,
       CAN_FIRE_RL_wsiS_ext_status_assign,
       CAN_FIRE_RL_wsiS_inc_tBusyCount,
       CAN_FIRE_RL_wsiS_operateD__dreg_update,
       CAN_FIRE_RL_wsiS_peerIsReady__dreg_update,
       CAN_FIRE_RL_wsiS_reqFifo__updateLevelCounter,
       CAN_FIRE_RL_wsiS_reqFifo_enq,
       CAN_FIRE_RL_wsiS_update_statusR,
       CAN_FIRE_RL_wsi_Es_doAlways,
       CAN_FIRE_RL_wsipass_doMessagePush,
       CAN_FIRE_wciS0_mAddr,
       CAN_FIRE_wciS0_mAddrSpace,
       CAN_FIRE_wciS0_mByteEn,
       CAN_FIRE_wciS0_mCmd,
       CAN_FIRE_wciS0_mData,
       CAN_FIRE_wciS0_mFlag,
       CAN_FIRE_wmemiM_sCmdAccept,
       CAN_FIRE_wmemiM_sData,
       CAN_FIRE_wmemiM_sDataAccept,
       CAN_FIRE_wmemiM_sResp,
       CAN_FIRE_wmemiM_sRespLast,
       CAN_FIRE_wsiM1_sReset_n,
       CAN_FIRE_wsiM1_sThreadBusy,
       CAN_FIRE_wsiS1_mBurstLength,
       CAN_FIRE_wsiS1_mBurstPrecise,
       CAN_FIRE_wsiS1_mByteEn,
       CAN_FIRE_wsiS1_mCmd,
       CAN_FIRE_wsiS1_mData,
       CAN_FIRE_wsiS1_mDataInfo,
       CAN_FIRE_wsiS1_mReqInfo,
       CAN_FIRE_wsiS1_mReqLast,
       CAN_FIRE_wsiS1_mReset_n,
       WILL_FIRE_RL_cycles_passed_count,
       WILL_FIRE_RL_delay_read_req,
       WILL_FIRE_RL_delay_read_resp,
       WILL_FIRE_RL_delay_write_req,
       WILL_FIRE_RL_delay_write_unblock,
       WILL_FIRE_RL_dlyReadCredit_accumulate,
       WILL_FIRE_RL_dlyWordsStored_accumulate,
       WILL_FIRE_RL_mesgRF_portA,
       WILL_FIRE_RL_mesgRF_portB,
       WILL_FIRE_RL_mesgRF_portB_read_data,
       WILL_FIRE_RL_mesgWF_portA,
       WILL_FIRE_RL_mesgWF_portB,
       WILL_FIRE_RL_mesgWF_portB_read_data,
       WILL_FIRE_RL_operating_actions,
       WILL_FIRE_RL_rdSer_begin,
       WILL_FIRE_RL_rdSer_body,
       WILL_FIRE_RL_rdSer_sync,
       WILL_FIRE_RL_wci_Es_doAlways_Req,
       WILL_FIRE_RL_wci_cfrd,
       WILL_FIRE_RL_wci_cfwr,
       WILL_FIRE_RL_wci_ctlAckReg__dreg_update,
       WILL_FIRE_RL_wci_ctl_op_complete,
       WILL_FIRE_RL_wci_ctl_op_start,
       WILL_FIRE_RL_wci_ctrl_EiI,
       WILL_FIRE_RL_wci_ctrl_IsO,
       WILL_FIRE_RL_wci_ctrl_OrE,
       WILL_FIRE_RL_wci_reqF__updateLevelCounter,
       WILL_FIRE_RL_wci_reqF_enq,
       WILL_FIRE_RL_wci_request_decode,
       WILL_FIRE_RL_wci_respF_both,
       WILL_FIRE_RL_wci_respF_decCtr,
       WILL_FIRE_RL_wci_respF_deq,
       WILL_FIRE_RL_wci_respF_incCtr,
       WILL_FIRE_RL_wci_sFlagReg__dreg_update,
       WILL_FIRE_RL_wci_sThreadBusy_reg,
       WILL_FIRE_RL_wmemi_Em_doAlways,
       WILL_FIRE_RL_wmemi_dhF_both,
       WILL_FIRE_RL_wmemi_dhF_decCtr,
       WILL_FIRE_RL_wmemi_dhF_deq,
       WILL_FIRE_RL_wmemi_dhF_incCtr,
       WILL_FIRE_RL_wmemi_operateD__dreg_update,
       WILL_FIRE_RL_wmemi_peerIsReady__dreg_update,
       WILL_FIRE_RL_wmemi_reqF_both,
       WILL_FIRE_RL_wmemi_reqF_decCtr,
       WILL_FIRE_RL_wmemi_reqF_deq,
       WILL_FIRE_RL_wmemi_reqF_incCtr,
       WILL_FIRE_RL_wmemi_respAdvance,
       WILL_FIRE_RL_wmemi_update_statusR,
       WILL_FIRE_RL_wmrd_mesgBegin,
       WILL_FIRE_RL_wmrd_mesgBodyResponse,
       WILL_FIRE_RL_wmwt_doAbort,
       WILL_FIRE_RL_wmwt_mesgBegin,
       WILL_FIRE_RL_wmwt_messageFinalize,
       WILL_FIRE_RL_wmwt_messagePushImprecise,
       WILL_FIRE_RL_wmwt_messagePushPrecise,
       WILL_FIRE_RL_wmwt_requestPrecise,
       WILL_FIRE_RL_wrtSer_begin,
       WILL_FIRE_RL_wrtSer_body,
       WILL_FIRE_RL_wsiM_ext_status_assign,
       WILL_FIRE_RL_wsiM_inc_tBusyCount,
       WILL_FIRE_RL_wsiM_operateD__dreg_update,
       WILL_FIRE_RL_wsiM_peerIsReady__dreg_update,
       WILL_FIRE_RL_wsiM_reqFifo_both,
       WILL_FIRE_RL_wsiM_reqFifo_decCtr,
       WILL_FIRE_RL_wsiM_reqFifo_deq,
       WILL_FIRE_RL_wsiM_reqFifo_incCtr,
       WILL_FIRE_RL_wsiM_sThreadBusy_reg,
       WILL_FIRE_RL_wsiM_update_statusR,
       WILL_FIRE_RL_wsiS_ext_status_assign,
       WILL_FIRE_RL_wsiS_inc_tBusyCount,
       WILL_FIRE_RL_wsiS_operateD__dreg_update,
       WILL_FIRE_RL_wsiS_peerIsReady__dreg_update,
       WILL_FIRE_RL_wsiS_reqFifo__updateLevelCounter,
       WILL_FIRE_RL_wsiS_reqFifo_enq,
       WILL_FIRE_RL_wsiS_update_statusR,
       WILL_FIRE_RL_wsi_Es_doAlways,
       WILL_FIRE_RL_wsipass_doMessagePush,
       WILL_FIRE_wciS0_mAddr,
       WILL_FIRE_wciS0_mAddrSpace,
       WILL_FIRE_wciS0_mByteEn,
       WILL_FIRE_wciS0_mCmd,
       WILL_FIRE_wciS0_mData,
       WILL_FIRE_wciS0_mFlag,
       WILL_FIRE_wmemiM_sCmdAccept,
       WILL_FIRE_wmemiM_sData,
       WILL_FIRE_wmemiM_sDataAccept,
       WILL_FIRE_wmemiM_sResp,
       WILL_FIRE_wmemiM_sRespLast,
       WILL_FIRE_wsiM1_sReset_n,
       WILL_FIRE_wsiM1_sThreadBusy,
       WILL_FIRE_wsiS1_mBurstLength,
       WILL_FIRE_wsiS1_mBurstPrecise,
       WILL_FIRE_wsiS1_mByteEn,
       WILL_FIRE_wsiS1_mCmd,
       WILL_FIRE_wsiS1_mData,
       WILL_FIRE_wsiS1_mDataInfo,
       WILL_FIRE_wsiS1_mReqInfo,
       WILL_FIRE_wsiS1_mReqLast,
       WILL_FIRE_wsiS1_mReset_n;

  // inputs to muxes for submodule ports
  reg [127 : 0] MUX_wide16Fa__enq_1__VAL_1, MUX_wide16Fa__enq_1__VAL_2;
  reg [33 : 0] MUX_wci_respF_q_0__write_1__VAL_2;
  wire [312 : 0] MUX_wsiM_reqFifo_q_0__write_1__VAL_1,
		 MUX_wsiM_reqFifo_q_0__write_1__VAL_2,
		 MUX_wsiM_reqFifo_q_1__write_1__VAL_1,
		 MUX_wsiM_reqFifo_x_wire__wset_1__VAL_1;
  wire [145 : 0] MUX_wmemi_dhF_q_0__write_1__VAL_1,
		 MUX_wmemi_dhF_q_0__write_1__VAL_2,
		 MUX_wmemi_dhF_q_1__write_1__VAL_1;
  wire [51 : 0] MUX_wmemi_reqF_q_0__write_1__VAL_1,
		MUX_wmemi_reqF_q_0__write_1__VAL_2,
		MUX_wmemi_reqF_q_1__write_1__VAL_1,
		MUX_wmemi_reqF_x_wire__wset_1__VAL_1,
		MUX_wmemi_reqF_x_wire__wset_1__VAL_2;
  wire [33 : 0] MUX_wci_respF_q_0__write_1__VAL_1,
		MUX_wci_respF_q_1__write_1__VAL_1,
		MUX_wci_respF_x_wire__wset_1__VAL_1,
		MUX_wci_respF_x_wire__wset_1__VAL_2;
  wire [31 : 0] MUX_mesgRdCount__write_1__VAL_1,
		MUX_mesgWtCount__write_1__VAL_1,
		MUX_metaWF__enq_1__VAL_1;
  wire [19 : 0] MUX_dlyRAG__write_1__VAL_1,
		MUX_dlyWAG__write_1__VAL_1,
		MUX_dlyWordsStored_value__write_1__VAL_2;
  wire [15 : 0] MUX_rdSerUnroll__write_1__VAL_2,
		MUX_unrollCnt__write_1__VAL_1,
		MUX_unrollCnt__write_1__VAL_2,
		MUX_wrtSerUnroll__write_1__VAL_1;
  wire [14 : 0] MUX_mesgLength__write_1__VAL_2, MUX_mesgLength__write_1__VAL_3;
  wire [13 : 0] MUX_mesgLengthSoFar__write_1__VAL_2;
  wire [11 : 0] MUX_wsiWordsRemain__write_1__VAL_2;
  wire [8 : 0] MUX_opcode__write_1__VAL_2;
  wire [7 : 0] MUX_dlyReadCredit_value__write_1__VAL_2;
  wire [1 : 0] MUX_rdSerPos__write_1__VAL_1,
	       MUX_wci_respF_c_r__write_1__VAL_1,
	       MUX_wci_respF_c_r__write_1__VAL_2,
	       MUX_wmemi_dhF_c_r__write_1__VAL_1,
	       MUX_wmemi_dhF_c_r__write_1__VAL_2,
	       MUX_wmemi_reqF_c_r__write_1__VAL_1,
	       MUX_wmemi_reqF_c_r__write_1__VAL_2,
	       MUX_wrtSerPos__write_1__VAL_1,
	       MUX_wrtSerPos__write_1__VAL_2,
	       MUX_wsiM_reqFifo_c_r__write_1__VAL_1,
	       MUX_wsiM_reqFifo_c_r__write_1__VAL_2;
  wire MUX_endOfMessage__write_1__SEL_1,
       MUX_impreciseBurst__write_1__SEL_2,
       MUX_mesgLength__write_1__SEL_2,
       MUX_mesgRdCount__write_1__SEL_1,
       MUX_metaWF__enq_1__SEL_1,
       MUX_rdSerEmpty__write_1__PSEL_1,
       MUX_rdSerEmpty__write_1__SEL_1,
       MUX_rdSyncWord__write_1__VAL_1,
       MUX_rdSyncWord__write_1__VAL_2,
       MUX_wci_illegalEdge__write_1__SEL_1,
       MUX_wci_illegalEdge__write_1__SEL_2,
       MUX_wci_illegalEdge__write_1__VAL_2,
       MUX_wci_respF_q_0__write_1__SEL_2,
       MUX_wci_respF_q_1__write_1__SEL_2,
       MUX_wide16Fa__enq_1__SEL_1,
       MUX_wmemi_dhF_q_0__write_1__SEL_2,
       MUX_wmemi_dhF_q_1__write_1__SEL_2,
       MUX_wmemi_reqF_q_0__write_1__SEL_2,
       MUX_wmemi_reqF_q_1__write_1__SEL_2,
       MUX_wrtSerStage__write_1__SEL_1,
       MUX_wrtSerStage_1__write_1__SEL_1,
       MUX_wrtSerStage_2__write_1__SEL_1,
       MUX_wrtSerStage_3__write_1__SEL_1,
       MUX_wsiM_reqFifo_q_0__write_1__SEL_2,
       MUX_wsiM_reqFifo_q_1__write_1__SEL_2;

  // remaining internal signals
  reg [63 : 0] v__h17561,
	       v__h17806,
	       v__h19118,
	       v__h19195,
	       v__h21672,
	       v__h2670,
	       v__h2817,
	       v__h3716;
  reg [31 : 0] x_data__h21804;
  reg CASE_wrtSerPos_0b1_0_1_1_1_2_1_3_0b1__q1,
      IF_wrtSerPos_11_EQ_0_12_OR_wrtSerPos_11_EQ_1_1_ETC___d904;
  wire [255 : 0] mesg__h22346, x__h15234, x__h16160, x__h19905;
  wire [127 : 0] IF_wrtSerPos_11_EQ_2_14_THEN_0x0_ELSE_mesgWF_w_ETC___d354,
		 IF_wrtSerPos_11_EQ_2_14_THEN_0x0_ELSE_metaWF_f_ETC___d377,
		 x1__h19969,
		 x1__h19978,
		 x1__h20492,
		 x1__h20501;
  wire [35 : 0] addr__h20994, addr__h21166;
  wire [31 : 0] rdat__h21847,
		rdat__h22030,
		rdat__h22038,
		rdat__h22046,
		rdat__h22054,
		v__h22720,
		x_byteEn__h22438;
  wire [23 : 0] x1_length__h17254, x__h21052, x__h21211, x__h21850;
  wire [13 : 0] mlp1__h17953, x__h17298;
  wire [11 : 0] x_burstLength__h22437;
  wire [10 : 0] x__h15126, x__h16052;
  wire [7 : 0] x1_opcode__h17253;
  wire [1 : 0] wrtSerPos_11_PLUS_1___d1014;
  wire NOT_dlyWordsStored_value_13_SLE_0_64_65_AND_NO_ETC___d272,
       NOT_mesgRF_rRdPtr_52_PLUS_512_93_EQ_mesgRF_rWr_ETC___d208,
       NOT_wsiS_reqFifo_countReg_96_ULE_1_97___d698,
       _dor1bytesWritten__EN_write,
       metaRF_RDY_enq__41_AND_NOT_rdSerEmpty_96_97_AN_ETC___d242,
       metaWF_RDY_deq__58_AND_NOT_wrtSerPos_11_EQ_3_1_ETC___d365,
       wci_cState_9_EQ_2_0_AND_dlyCtrl_4_BITS_3_TO_0__ETC___d397;

  // action method wciS0_mCmd
  assign CAN_FIRE_wciS0_mCmd = 1'b1 ;
  assign WILL_FIRE_wciS0_mCmd = 1'b1 ;

  // action method wciS0_mAddrSpace
  assign CAN_FIRE_wciS0_mAddrSpace = 1'b1 ;
  assign WILL_FIRE_wciS0_mAddrSpace = 1'b1 ;

  // action method wciS0_mByteEn
  assign CAN_FIRE_wciS0_mByteEn = 1'b1 ;
  assign WILL_FIRE_wciS0_mByteEn = 1'b1 ;

  // action method wciS0_mAddr
  assign CAN_FIRE_wciS0_mAddr = 1'b1 ;
  assign WILL_FIRE_wciS0_mAddr = 1'b1 ;

  // action method wciS0_mData
  assign CAN_FIRE_wciS0_mData = 1'b1 ;
  assign WILL_FIRE_wciS0_mData = 1'b1 ;

  // value method wciS0_sResp
  assign wciS0_SResp = wci_respF_q_0[33:32] ;

  // value method wciS0_sData
  assign wciS0_SData = wci_respF_q_0[31:0] ;

  // value method wciS0_sThreadBusy
  assign wciS0_SThreadBusy = wci_reqF_countReg > 2'b01 || wci_isReset__VAL ;

  // value method wciS0_sFlag
  assign wciS0_SFlag = { 1'b1, wci_sFlagReg } ;

  // action method wciS0_mFlag
  assign CAN_FIRE_wciS0_mFlag = 1'b1 ;
  assign WILL_FIRE_wciS0_mFlag = 1'b1 ;

  // action method wsiS1_mCmd
  assign CAN_FIRE_wsiS1_mCmd = 1'b1 ;
  assign WILL_FIRE_wsiS1_mCmd = 1'b1 ;

  // action method wsiS1_mReqLast
  assign CAN_FIRE_wsiS1_mReqLast = 1'b1 ;
  assign WILL_FIRE_wsiS1_mReqLast = wsiS1_MReqLast ;

  // action method wsiS1_mBurstPrecise
  assign CAN_FIRE_wsiS1_mBurstPrecise = 1'b1 ;
  assign WILL_FIRE_wsiS1_mBurstPrecise = wsiS1_MBurstPrecise ;

  // action method wsiS1_mBurstLength
  assign CAN_FIRE_wsiS1_mBurstLength = 1'b1 ;
  assign WILL_FIRE_wsiS1_mBurstLength = 1'b1 ;

  // action method wsiS1_mData
  assign CAN_FIRE_wsiS1_mData = 1'b1 ;
  assign WILL_FIRE_wsiS1_mData = 1'b1 ;

  // action method wsiS1_mByteEn
  assign CAN_FIRE_wsiS1_mByteEn = 1'b1 ;
  assign WILL_FIRE_wsiS1_mByteEn = 1'b1 ;

  // action method wsiS1_mReqInfo
  assign CAN_FIRE_wsiS1_mReqInfo = 1'b1 ;
  assign WILL_FIRE_wsiS1_mReqInfo = 1'b1 ;

  // action method wsiS1_mDataInfo
  assign CAN_FIRE_wsiS1_mDataInfo = 1'b1 ;
  assign WILL_FIRE_wsiS1_mDataInfo = 1'b1 ;

  // value method wsiS1_sThreadBusy
  assign wsiS1_SThreadBusy =
	     NOT_wsiS_reqFifo_countReg_96_ULE_1_97___d698 ||
	     wsiS_isReset__VAL ||
	     !wsiS_operateD ||
	     !wsiS_peerIsReady ;

  // value method wsiS1_sReset_n
  assign wsiS1_SReset_n = !wsiS_isReset__VAL && wsiS_operateD ;

  // action method wsiS1_mReset_n
  assign CAN_FIRE_wsiS1_mReset_n = 1'b1 ;
  assign WILL_FIRE_wsiS1_mReset_n = wsiS1_MReset_n ;

  // value method wsiM1_mCmd
  assign wsiM1_MCmd = wsiM_sThreadBusy_d ? 3'b000 : wsiM_reqFifo_q_0[312:310] ;

  // value method wsiM1_mReqLast
  assign wsiM1_MReqLast = !wsiM_sThreadBusy_d && wsiM_reqFifo_q_0[309] ;

  // value method wsiM1_mBurstPrecise
  assign wsiM1_MBurstPrecise = !wsiM_sThreadBusy_d && wsiM_reqFifo_q_0[308] ;

  // value method wsiM1_mBurstLength
  assign wsiM1_MBurstLength =
	     wsiM_sThreadBusy_d ? 12'b00 : wsiM_reqFifo_q_0[307:296] ;

  // value method wsiM1_mData
  assign wsiM1_MData = wsiM_reqFifo_q_0[295:40] ;

  // value method wsiM1_mByteEn
  assign wsiM1_MByteEn = wsiM_reqFifo_q_0[39:8] ;

  // value method wsiM1_mReqInfo
  assign wsiM1_MReqInfo = wsiM_sThreadBusy_d ? 8'b00000000 : wsiM_reqFifo_q_0[7:0] ;

  // action method wsiM1_sThreadBusy
  assign CAN_FIRE_wsiM1_sThreadBusy = 1'b1 ;
  assign WILL_FIRE_wsiM1_sThreadBusy = wsiM1_SThreadBusy ;

  // value method wsiM1_mReset_n
  assign wsiM1_MReset_n = !wsiM_isReset__VAL && wsiM_operateD ;

  // action method wsiM1_sReset_n
  assign CAN_FIRE_wsiM1_sReset_n = 1'b1 ;
  assign WILL_FIRE_wsiM1_sReset_n = wsiM1_SReset_n ;

  // value method wmemiM_mCmd
  assign wmemiM_MCmd = wmemi_reqF_q_0[51:49] ;

  // value method wmemiM_mReqLast
  assign wmemiM_MReqLast = wmemi_reqF_q_0[48] ;

  // value method wmemiM_mAddr
  assign wmemiM_MAddr = wmemi_reqF_q_0[47:12] ;

  // value method wmemiM_mBurstLength
  assign wmemiM_MBurstLength = wmemi_reqF_q_0[11:0] ;

  // value method wmemiM_mDataValid
  assign wmemiM_MDataValid = wmemi_dhF_q_0[145] ;

  // value method wmemiM_mDataLast
  assign wmemiM_MDataLast = wmemi_dhF_q_0[144] ;

  // value method wmemiM_mData
  assign wmemiM_MData = wmemi_dhF_q_0[143:16] ;

  // value method wmemiM_mDataByteEn
  assign wmemiM_MDataByteEn = wmemi_dhF_q_0[15:0] ;

  // action method wmemiM_sResp
  assign CAN_FIRE_wmemiM_sResp = 1'b1 ;
  assign WILL_FIRE_wmemiM_sResp = 1'b1 ;

  // action method wmemiM_sRespLast
  assign CAN_FIRE_wmemiM_sRespLast = 1'b1 ;
  assign WILL_FIRE_wmemiM_sRespLast = wmemiM_SRespLast ;

  // action method wmemiM_sData
  assign CAN_FIRE_wmemiM_sData = 1'b1 ;
  assign WILL_FIRE_wmemiM_sData = 1'b1 ;

  // action method wmemiM_sCmdAccept
  assign CAN_FIRE_wmemiM_sCmdAccept = 1'b1 ;
  assign WILL_FIRE_wmemiM_sCmdAccept = wmemiM_SCmdAccept ;

  // action method wmemiM_sDataAccept
  assign CAN_FIRE_wmemiM_sDataAccept = 1'b1 ;
  assign WILL_FIRE_wmemiM_sDataAccept = wmemiM_SDataAccept ;

  // value method wmemiM_mReset_n
  assign wmemiM_MReset_n = !wmemi_isReset__VAL && wmemi_operateD ;

  // submodule mesgRF_memory
  
// #(.PIPELINED(1'b0),
//	  .ADDR_WIDTH(32'b010),
//	  .DATA_WIDTH(32'b1056),
//	  .MEMSIZE(11'b1024)) mesgRF_memory

wire [255:0] dp_out_not_used1;
wire [255:0] dp_out_not_used2;

  dual_port_ram #( .ADDR_WIDTH(10), .DATA_WIDTH(256)) dpram1 (
        					.clk(wciS0_Clk),
        				    .addr1(mesgRF_memory__ADDRA),
        				    .addr2(mesgRF_memory__ADDRB),
        				    .data1(mesgRF_memory__DIA),
        				    .data2(mesgRF_memory__DIB),
        				    .we1(mesgRF_memory__WEA),
        				    .we2(mesgRF_memory__WEB),
        				    .out1(dp_out_not_used1),
        				    .out2(mesgRF_memory__DOB)
        					);

  // submodule mesgWF_memory
//#(.PIPELINED(1'b0),
//	  .ADDR_WIDTH(32'b010),
//	  .DATA_WIDTH(32'b1056),
//	  .MEMSIZE(11'b1024)) mesgWF_memory(
	  
 dual_port_ram #( .ADDR_WIDTH(10), .DATA_WIDTH(256)) dpram2   (
        					.clk(wciS0_Clk),
        				    .addr1(mesgWF_memory__ADDRA),
        				    .addr2(mesgWF_memory__ADDRB),
        				    .data1(mesgWF_memory__DIA),
        				    .data2(mesgWF_memory__DIB),
        				    .we1(mesgWF_memory__WEA),
        				    .we2(mesgWF_memory__WEB),
        				    .out1(dp_out_not_used2),
        				    .out2(mesgWF_memory__DOB)
        					);

  // submodule metaRF
  arSRLFIFO_a 	ars1	(
					 .CLK(wciS0_Clk),
				     .RST_N(wciS0_MReset_n),
				     .D_IN(metaRF__D_IN),
				     .ENQ(metaRF__ENQ),
				     .DEQ(metaRF__DEQ),
				     .CLR(metaRF__CLR),
				     .D_OUT(metaRF__D_OUT),
				     .EMPTY_N(metaRF__EMPTY_N),
				     .FULL_N(metaRF__FULL_N)
					 );

  // submodule metaWF
  arSRLFIFO_b 	ars2	(
					 .CLK(wciS0_Clk),
				     .RST_N(wciS0_MReset_n),
				     .D_IN(metaWF__D_IN),
				     .ENQ(metaWF__ENQ),
				     .DEQ(metaWF__DEQ),
				     .CLR(metaWF__CLR),
				     .D_OUT(metaWF__D_OUT),
				     .EMPTY_N(metaWF__EMPTY_N),
				     .FULL_N(metaWF__FULL_N)
					 );

  // submodule wci_isReset
  ResetToBool wci_isReset(.RST(wciS0_MReset_n), .VAL(wci_isReset__VAL));

  wire full_a_not_used;
  // submodule wci_reqF
  SizedFIFO_a 	sizefifo1	(
					.CLK(wciS0_Clk),
					.D_IN(wci_reqF__D_IN),
					.ENQ(wci_reqF__ENQ),
					.DEQ(wci_reqF__DEQ),
					.CLR(wci_reqF__CLR),
					.D_OUT(wci_reqF__D_OUT),
					.FULL_N(full_a_not_used),
					.EMPTY_N(wci_reqF__EMPTY_N)
					);

  // submodule wide16Fa
  arSRLFIFO_c ars3		(
						.CLK(wciS0_Clk),
				       .RST_N(wciS0_MReset_n),
				       .D_IN(wide16Fa__D_IN),
				       .ENQ(wide16Fa__ENQ),
				       .DEQ(wide16Fa__DEQ),
				       .CLR(wide16Fa__CLR),
				       .D_OUT(wide16Fa__D_OUT),
				       .EMPTY_N(wide16Fa__EMPTY_N),
				       .FULL_N(wide16Fa__FULL_N)
					   );

  // submodule wide16Fb
  arSRLFIFO_d ars4		(
						.CLK(wciS0_Clk),
				       .RST_N(wciS0_MReset_n),
				       .D_IN(wide16Fb__D_IN),
				       .ENQ(wide16Fb__ENQ),
				       .DEQ(wide16Fb__DEQ),
				       .CLR(wide16Fb__CLR),
				       .D_OUT(wide16Fb__D_OUT),
				       .EMPTY_N(wide16Fb__EMPTY_N),
				       .FULL_N(wide16Fb__FULL_N)
					   );

  // submodule wmemi_isReset
  ResetToBool wmemi_isReset(.RST(wciS0_MReset_n), .VAL(wmemi_isReset__VAL));

  // submodule wmemi_respF
//   #(.width(32'b0131),
//	  .guarded(32'b01)) wmemi_respF(.RST_N(wciS0_MReset_n),
  SizedFIFO_x	fifo_2		(
				       .CLK(wciS0_Clk),
				       .D_IN(wmemi_respF__D_IN),
				       .ENQ(wmemi_respF__ENQ),
				       .DEQ(wmemi_respF__DEQ),
				       .CLR(wmemi_respF__CLR),
				       .D_OUT(wmemi_respF__D_OUT),
				       .FULL_N(wmemi_respF__FULL_N),
				       .EMPTY_N(wmemi_respF__EMPTY_N)
					   );

  // submodule wsiM_isReset
  ResetToBool wsiM_isReset(.RST(wciS0_MReset_n), .VAL(wsiM_isReset__VAL));

  // submodule wsiS_isReset
  ResetToBool wsiS_isReset(.RST(wciS0_MReset_n), .VAL(wsiS_isReset__VAL));

  //#(.p1width(32'b1113),
	//      .p2depth(32'b11),
	//      .p3cntr_width(32'b01),
	//      .guarded(32'b01)) wsiS_reqFifo(.RST_N(wciS0_MReset_n),
  // submodule wsiS_reqFifo
  SizedFIFO_b sizefifo2 (
						.CLK(wciS0_Clk),
					    .D_IN(wsiS_reqFifo__D_IN),
					    .ENQ(wsiS_reqFifo__ENQ),
					    .DEQ(wsiS_reqFifo__DEQ),
					    .CLR(wsiS_reqFifo__CLR),
					    .D_OUT(wsiS_reqFifo__D_OUT),
					    .FULL_N(wsiS_reqFifo__FULL_N),
					    .EMPTY_N(wsiS_reqFifo__EMPTY_N)
						);

  // rule RL_wci_request_decode
  assign CAN_FIRE_RL_wci_request_decode = wci_reqF__EMPTY_N ;
  assign WILL_FIRE_RL_wci_request_decode = wci_reqF__EMPTY_N ;

  // rule RL_wci_ctl_op_start
  assign CAN_FIRE_RL_wci_ctl_op_start =
	     wci_reqF__EMPTY_N && wci_wci_ctrl_pw__whas ;
  assign WILL_FIRE_RL_wci_ctl_op_start =
	     CAN_FIRE_RL_wci_ctl_op_start &&
	     !WILL_FIRE_RL_wci_ctl_op_complete ;

  // rule RL_wci_ctrl_EiI
  assign CAN_FIRE_RL_wci_ctrl_EiI =
	     wci_wci_ctrl_pw__whas && WILL_FIRE_RL_wci_ctl_op_start &&
	     wci_cState == 3'b000 &&
	     wci_reqF__D_OUT[36:34] == 3'b000 ;
  assign WILL_FIRE_RL_wci_ctrl_EiI = CAN_FIRE_RL_wci_ctrl_EiI ;

  // rule RL_wci_ctrl_OrE
  assign CAN_FIRE_RL_wci_ctrl_OrE =
	     wci_wci_ctrl_pw__whas && WILL_FIRE_RL_wci_ctl_op_start &&
	     wci_cState == 3'b010 &&
	     wci_reqF__D_OUT[36:34] == 3'b011 ;
  assign WILL_FIRE_RL_wci_ctrl_OrE = CAN_FIRE_RL_wci_ctrl_OrE ;

  // rule RL_wci_respF_deq
  assign CAN_FIRE_RL_wci_respF_deq = 1'b1 ;
  assign WILL_FIRE_RL_wci_respF_deq = 1'b1 ;

  // rule RL_wmemi_update_statusR
  assign CAN_FIRE_RL_wmemi_update_statusR = 1'b1 ;
  assign WILL_FIRE_RL_wmemi_update_statusR = 1'b1 ;

  // rule RL_wci_sThreadBusy_reg
  assign CAN_FIRE_RL_wci_sThreadBusy_reg = 1'b1 ;
  assign WILL_FIRE_RL_wci_sThreadBusy_reg = 1'b1 ;

  // rule RL_wci_sFlagReg__dreg_update
  assign CAN_FIRE_RL_wci_sFlagReg__dreg_update = 1'b1 ;
  assign WILL_FIRE_RL_wci_sFlagReg__dreg_update = 1'b1 ;

  // rule RL_wsi_Es_doAlways
  assign CAN_FIRE_RL_wsi_Es_doAlways = 1'b1 ;
  assign WILL_FIRE_RL_wsi_Es_doAlways = 1'b1 ;

  // rule RL_wsiS_update_statusR
  assign CAN_FIRE_RL_wsiS_update_statusR = 1'b1 ;
  assign WILL_FIRE_RL_wsiS_update_statusR = 1'b1 ;

  // rule RL_wsiS_ext_status_assign
  assign CAN_FIRE_RL_wsiS_ext_status_assign = 1'b1 ;
  assign WILL_FIRE_RL_wsiS_ext_status_assign = 1'b1 ;

  // rule RL_wsiS_inc_tBusyCount
  assign CAN_FIRE_RL_wsiS_inc_tBusyCount =
	     wsiS_operateD && wsiS_peerIsReady &&
	     NOT_wsiS_reqFifo_countReg_96_ULE_1_97___d698 ;
  assign WILL_FIRE_RL_wsiS_inc_tBusyCount = CAN_FIRE_RL_wsiS_inc_tBusyCount ;

  // rule RL_wsiS_reqFifo_enq
  assign CAN_FIRE_RL_wsiS_reqFifo_enq =
	     wsiS_operateD && wsiS_peerIsReady &&
	     wsiS_wsiReq__wget[312:310] == 3'b001 ;
  assign WILL_FIRE_RL_wsiS_reqFifo_enq = CAN_FIRE_RL_wsiS_reqFifo_enq ;

  // rule RL_wsiS_peerIsReady__dreg_update
  assign CAN_FIRE_RL_wsiS_peerIsReady__dreg_update = 1'b1 ;
  assign WILL_FIRE_RL_wsiS_peerIsReady__dreg_update = 1'b1 ;

  // rule RL_wsiM_update_statusR
  assign CAN_FIRE_RL_wsiM_update_statusR = 1'b1 ;
  assign WILL_FIRE_RL_wsiM_update_statusR = 1'b1 ;

  // rule RL_wsiM_ext_status_assign
  assign CAN_FIRE_RL_wsiM_ext_status_assign = 1'b1 ;
  assign WILL_FIRE_RL_wsiM_ext_status_assign = 1'b1 ;

  // rule RL_wci_cfrd
  assign CAN_FIRE_RL_wci_cfrd =
	     wci_respF_c_r != 2'b10 && wci_reqF__EMPTY_N &&
	     wci_wci_cfrd_pw__whas ;
  assign WILL_FIRE_RL_wci_cfrd =
	     CAN_FIRE_RL_wci_cfrd && !WILL_FIRE_RL_wci_ctl_op_start &&
	     !WILL_FIRE_RL_wci_ctl_op_complete ;

  // rule RL_wsiM_inc_tBusyCount
  assign CAN_FIRE_RL_wsiM_inc_tBusyCount =
	     wsiM_operateD && wsiM_peerIsReady && wsiM_sThreadBusy_d ;
  assign WILL_FIRE_RL_wsiM_inc_tBusyCount = CAN_FIRE_RL_wsiM_inc_tBusyCount ;

  // rule RL_wsiM_reqFifo_deq
  assign CAN_FIRE_RL_wsiM_reqFifo_deq =
	     wsiM_reqFifo_c_r != 2'b00 && !wsiM_sThreadBusy_d ;
  assign WILL_FIRE_RL_wsiM_reqFifo_deq = CAN_FIRE_RL_wsiM_reqFifo_deq ;

  // rule RL_wsiM_sThreadBusy_reg
  assign CAN_FIRE_RL_wsiM_sThreadBusy_reg = 1'b1 ;
  assign WILL_FIRE_RL_wsiM_sThreadBusy_reg = 1'b1 ;

  // rule RL_wsiM_peerIsReady__dreg_update
  assign CAN_FIRE_RL_wsiM_peerIsReady__dreg_update = 1'b1 ;
  assign WILL_FIRE_RL_wsiM_peerIsReady__dreg_update = 1'b1 ;

  // rule RL_operating_actions
  assign CAN_FIRE_RL_operating_actions = wci_cState == 3'b010 ;
  assign WILL_FIRE_RL_operating_actions = wci_cState == 3'b010 ;

  // rule RL_wsiS_operateD__dreg_update
  assign CAN_FIRE_RL_wsiS_operateD__dreg_update = 1'b1 ;
  assign WILL_FIRE_RL_wsiS_operateD__dreg_update = 1'b1 ;

  // rule RL_wsiM_operateD__dreg_update
  assign CAN_FIRE_RL_wsiM_operateD__dreg_update = 1'b1 ;
  assign WILL_FIRE_RL_wsiM_operateD__dreg_update = 1'b1 ;

  // rule RL_wmrd_mesgBegin
  assign CAN_FIRE_RL_wmrd_mesgBegin =
	     metaRF__EMPTY_N && wci_cState == 3'b010 && dlyCtrl[3:0] == 4'h7 &&
	     unrollCnt == 16'b0000000000000000 ;
  assign WILL_FIRE_RL_wmrd_mesgBegin = CAN_FIRE_RL_wmrd_mesgBegin ;

  // rule RL_wmwt_messageFinalize
  assign CAN_FIRE_RL_wmwt_messageFinalize =
	     (!impreciseBurst || metaWF__FULL_N) &&
	     wci_cState_9_EQ_2_0_AND_dlyCtrl_4_BITS_3_TO_0__ETC___d397 ;
  assign WILL_FIRE_RL_wmwt_messageFinalize =
	     CAN_FIRE_RL_wmwt_messageFinalize ;

  // rule RL_wci_Es_doAlways_Req
  assign CAN_FIRE_RL_wci_Es_doAlways_Req = 1'b1 ;
  assign WILL_FIRE_RL_wci_Es_doAlways_Req = 1'b1 ;

  // rule RL_wci_reqF_enq
  assign CAN_FIRE_RL_wci_reqF_enq = wci_wciReq__wget[59:57] != 3'b000 ;
  assign WILL_FIRE_RL_wci_reqF_enq = CAN_FIRE_RL_wci_reqF_enq ;

  // rule RL_wsipass_doMessagePush
  assign CAN_FIRE_RL_wsipass_doMessagePush =
	     wsiM_reqFifo_c_r != 2'b10 && wsiS_reqFifo__EMPTY_N &&
	     wci_cState == 3'b010 &&
	     dlyCtrl[3:0] == 4'h0 ;
  assign WILL_FIRE_RL_wsipass_doMessagePush =
	     CAN_FIRE_RL_wsipass_doMessagePush ;

  // rule RL_delay_write_req
  assign CAN_FIRE_RL_delay_write_req =
	     wide16Fa__EMPTY_N && wmemi_reqF_c_r != 2'b10 &&
	     wmemi_dhF_c_r != 2'b10 &&
	     wmemi_operateD &&
	     wmemi_peerIsReady &&
	     wci_cState == 3'b010 &&
	     dlyCtrl[3:0] == 4'h7 &&
	     !blockDelayWrite ;
  assign WILL_FIRE_RL_delay_write_req = CAN_FIRE_RL_delay_write_req ;

  // rule RL_delay_read_req
  assign CAN_FIRE_RL_delay_read_req =
	     wmemi_reqF_c_r != 2'b10 && wmemi_operateD && wmemi_peerIsReady &&
	     wci_cState == 3'b010 &&
	     dlyCtrl[3:0] == 4'h7 &&
	     NOT_dlyWordsStored_value_13_SLE_0_64_65_AND_NO_ETC___d272 &&
	     (dlyReadCredit_value ^ 8'h80) > 8'b10000000 ;
  assign WILL_FIRE_RL_delay_read_req =
	     CAN_FIRE_RL_delay_read_req && !WILL_FIRE_RL_delay_write_req ;

  // rule RL_wmwt_messagePushPrecise
  assign CAN_FIRE_RL_wmwt_messagePushPrecise =
	     mesgWF_rRdPtr + 11'b01000000000 != mesgWF_rWrPtr &&
	     wsiS_reqFifo__EMPTY_N &&
	     wci_cState == 3'b010 &&
	     dlyCtrl[3:0] == 4'h7 &&
	     wsiWordsRemain != 12'b00 &&
	     mesgReqValid &&
	     preciseBurst ;
  assign WILL_FIRE_RL_wmwt_messagePushPrecise =
	     CAN_FIRE_RL_wmwt_messagePushPrecise &&
	     !WILL_FIRE_RL_wmwt_messagePushImprecise &&
	     !WILL_FIRE_RL_wmwt_messageFinalize ;

  // rule RL_wmwt_requestPrecise
  assign CAN_FIRE_RL_wmwt_requestPrecise =
	     metaWF__FULL_N && wci_cState == 3'b010 && dlyCtrl[3:0] == 4'h7 &&
	     readyToRequest &&
	     preciseBurst ;
  assign WILL_FIRE_RL_wmwt_requestPrecise =
	     CAN_FIRE_RL_wmwt_requestPrecise &&
	     !WILL_FIRE_RL_wmwt_messageFinalize ;

  // rule RL_wmwt_messagePushImprecise
  assign CAN_FIRE_RL_wmwt_messagePushImprecise =
	     mesgWF_rRdPtr + 11'b01000000000 != mesgWF_rWrPtr &&
	     wsiS_reqFifo__EMPTY_N &&
	     wci_cState == 3'b010 &&
	     dlyCtrl[3:0] == 4'h7 &&
	     readyToPush &&
	     impreciseBurst ;
  assign WILL_FIRE_RL_wmwt_messagePushImprecise =
	     CAN_FIRE_RL_wmwt_messagePushImprecise &&
	     !WILL_FIRE_RL_wmwt_messageFinalize ;

  // rule RL_wsiS_reqFifo__updateLevelCounter
  assign CAN_FIRE_RL_wsiS_reqFifo__updateLevelCounter =
	     CAN_FIRE_RL_wsiS_reqFifo_enq != wsiS_reqFifo_r_deq__whas ;
  assign WILL_FIRE_RL_wsiS_reqFifo__updateLevelCounter =
	     CAN_FIRE_RL_wsiS_reqFifo__updateLevelCounter ;

  // rule RL_wmwt_mesgBegin
  assign CAN_FIRE_RL_wmwt_mesgBegin =
	     wsiS_reqFifo__EMPTY_N && wci_cState == 3'b010 &&
	     dlyCtrl[3:0] == 4'h7 &&
	     !opcode[8] ;
  assign WILL_FIRE_RL_wmwt_mesgBegin =
	     CAN_FIRE_RL_wmwt_mesgBegin &&
	     !WILL_FIRE_RL_wmwt_messagePushPrecise &&
	     !WILL_FIRE_RL_wmwt_messagePushImprecise &&
	     !WILL_FIRE_RL_wmwt_messageFinalize ;

  // rule RL_wmwt_doAbort
  assign CAN_FIRE_RL_wmwt_doAbort =
	     wci_cState == 3'b010 && dlyCtrl[3:0] == 4'h7 && doAbort ;
  assign WILL_FIRE_RL_wmwt_doAbort = CAN_FIRE_RL_wmwt_doAbort ;

  // rule RL_wmemi_Em_doAlways
  assign CAN_FIRE_RL_wmemi_Em_doAlways = 1'b1 ;
  assign WILL_FIRE_RL_wmemi_Em_doAlways = 1'b1 ;

  // rule RL_rdSer_sync
  assign CAN_FIRE_RL_rdSer_sync =
	     wci_cState == 3'b010 && dlyCtrl[3:0] == 4'h7 && rdSyncWord ;
  assign WILL_FIRE_RL_rdSer_sync = CAN_FIRE_RL_rdSer_sync ;

  // rule RL_rdSer_body
  assign CAN_FIRE_RL_rdSer_body =
	     NOT_mesgRF_rRdPtr_52_PLUS_512_93_EQ_mesgRF_rWr_ETC___d208 &&
	     wci_cState == 3'b010 &&
	     dlyCtrl[3:0] == 4'h7 &&
	     rdSerUnroll != 16'b0000000000000000 &&
	     !rdSyncWord ;
  assign WILL_FIRE_RL_rdSer_body = CAN_FIRE_RL_rdSer_body ;

  // rule RL_rdSer_begin
  assign CAN_FIRE_RL_rdSer_begin =
	     metaRF_RDY_enq__41_AND_NOT_rdSerEmpty_96_97_AN_ETC___d242 &&
	     wci_cState == 3'b010 &&
	     dlyCtrl[3:0] == 4'h7 &&
	     rdSerUnroll == 16'b0000000000000000 &&
	     !rdSyncWord ;
  assign WILL_FIRE_RL_rdSer_begin = CAN_FIRE_RL_rdSer_begin ;

  // rule RL_delay_read_resp
  assign CAN_FIRE_RL_delay_read_resp =
	     wide16Fb__FULL_N && wmemi_respF__EMPTY_N && wci_cState == 3'b010 &&
	     dlyCtrl[3:0] == 4'h7 ;
  assign WILL_FIRE_RL_delay_read_resp = CAN_FIRE_RL_delay_read_resp ;

  // rule RL_delay_write_unblock
  assign CAN_FIRE_RL_delay_write_unblock =
	     wci_cState == 3'b010 && dlyCtrl[3:0] == 4'h7 && blockDelayWrite ;
  assign WILL_FIRE_RL_delay_write_unblock = CAN_FIRE_RL_delay_write_unblock ;

  // rule RL_wrtSer_begin
  assign CAN_FIRE_RL_wrtSer_begin =
	     metaWF__EMPTY_N &&
	     metaWF_RDY_deq__58_AND_NOT_wrtSerPos_11_EQ_3_1_ETC___d365 &&
	     wci_cState == 3'b010 &&
	     dlyCtrl[3:0] == 4'h7 &&
	     wrtSerUnroll == 16'b0000000000000000 ;
  assign WILL_FIRE_RL_wrtSer_begin = CAN_FIRE_RL_wrtSer_begin ;

  // rule RL_cycles_passed_count
  assign CAN_FIRE_RL_cycles_passed_count = wsiS_statusR[0] ;
  assign WILL_FIRE_RL_cycles_passed_count = CAN_FIRE_RL_cycles_passed_count ;

  // rule RL_dlyWordsStored_accumulate
  assign CAN_FIRE_RL_dlyWordsStored_accumulate = 1'b1 ;
  assign WILL_FIRE_RL_dlyWordsStored_accumulate = 1'b1 ;

  // rule RL_dlyReadCredit_accumulate
  assign CAN_FIRE_RL_dlyReadCredit_accumulate = 1'b1 ;
  assign WILL_FIRE_RL_dlyReadCredit_accumulate = 1'b1 ;

  // rule RL_wci_ctrl_IsO
  assign CAN_FIRE_RL_wci_ctrl_IsO =
	     wci_wci_ctrl_pw__whas && WILL_FIRE_RL_wci_ctl_op_start &&
	     wci_cState == 3'b001 &&
	     wci_reqF__D_OUT[36:34] == 3'b001 ;
  assign WILL_FIRE_RL_wci_ctrl_IsO = CAN_FIRE_RL_wci_ctrl_IsO ;

  // rule RL_mesgRF_portB_read_data
  assign CAN_FIRE_RL_mesgRF_portB_read_data = 1'b1 ;
  assign WILL_FIRE_RL_mesgRF_portB_read_data = 1'b1 ;

  // rule RL_wmrd_mesgBodyResponse
  assign CAN_FIRE_RL_wmrd_mesgBodyResponse =
	     wsiM_reqFifo_c_r != 2'b10 && mesgRF_rRdPtr != mesgRF_rWrPtr &&
	     wci_cState == 3'b010 &&
	     dlyCtrl[3:0] == 4'h7 &&
	     unrollCnt != 16'b0000000000000000 ;
  assign WILL_FIRE_RL_wmrd_mesgBodyResponse =
	     CAN_FIRE_RL_wmrd_mesgBodyResponse ;

  // rule RL_wsiM_reqFifo_both
  assign CAN_FIRE_RL_wsiM_reqFifo_both =
	     ((wsiM_reqFifo_c_r == 2'b01) ?
		wsiM_reqFifo_x_wire__whas :
		wsiM_reqFifo_c_r != 2'b10 || wsiM_reqFifo_x_wire__whas) &&
	     CAN_FIRE_RL_wsiM_reqFifo_deq &&
	     wsiM_reqFifo_enqueueing__whas ;
  assign WILL_FIRE_RL_wsiM_reqFifo_both = CAN_FIRE_RL_wsiM_reqFifo_both ;

  // rule RL_wsiM_reqFifo_decCtr
  assign CAN_FIRE_RL_wsiM_reqFifo_decCtr =
	     CAN_FIRE_RL_wsiM_reqFifo_deq && !wsiM_reqFifo_enqueueing__whas ;
  assign WILL_FIRE_RL_wsiM_reqFifo_decCtr = CAN_FIRE_RL_wsiM_reqFifo_decCtr ;

  // rule RL_wsiM_reqFifo_incCtr
  assign CAN_FIRE_RL_wsiM_reqFifo_incCtr =
	     ((wsiM_reqFifo_c_r == 2'b00) ?
		wsiM_reqFifo_x_wire__whas :
		wsiM_reqFifo_c_r != 2'b01 || wsiM_reqFifo_x_wire__whas) &&
	     wsiM_reqFifo_enqueueing__whas &&
	     !CAN_FIRE_RL_wsiM_reqFifo_deq ;
  assign WILL_FIRE_RL_wsiM_reqFifo_incCtr = CAN_FIRE_RL_wsiM_reqFifo_incCtr ;

  // rule RL_mesgRF_portB
  assign CAN_FIRE_RL_mesgRF_portB = 1'b1 ;
  assign WILL_FIRE_RL_mesgRF_portB = 1'b1 ;

  // rule RL_mesgRF_portA
  assign CAN_FIRE_RL_mesgRF_portA = 1'b1 ;
  assign WILL_FIRE_RL_mesgRF_portA = 1'b1 ;

  // rule RL_mesgWF_portB_read_data
  assign CAN_FIRE_RL_mesgWF_portB_read_data = 1'b1 ;
  assign WILL_FIRE_RL_mesgWF_portB_read_data = 1'b1 ;

  // rule RL_wrtSer_body
  assign CAN_FIRE_RL_wrtSer_body =
	     mesgWF_rRdPtr != mesgWF_rWrPtr &&
	     CASE_wrtSerPos_0b1_0_1_1_1_2_1_3_0b1__q1 &&
	     (wrtSerPos != 2'b11 && wrtSerUnroll != 16'b0000000000000001 ||
	      IF_wrtSerPos_11_EQ_0_12_OR_wrtSerPos_11_EQ_1_1_ETC___d904) &&
	     wci_cState == 3'b010 &&
	     dlyCtrl[3:0] == 4'h7 &&
	     wrtSerUnroll != 16'b0000000000000000 ;
  assign WILL_FIRE_RL_wrtSer_body = CAN_FIRE_RL_wrtSer_body ;

  // rule RL_wci_ctl_op_complete
  assign CAN_FIRE_RL_wci_ctl_op_complete =
	     wci_respF_c_r != 2'b10 && wci_ctlOpActive && wci_ctlAckReg ;
  assign WILL_FIRE_RL_wci_ctl_op_complete = CAN_FIRE_RL_wci_ctl_op_complete ;

  // rule RL_wci_cfwr
  assign CAN_FIRE_RL_wci_cfwr =
	     wci_respF_c_r != 2'b10 && wci_reqF__EMPTY_N &&
	     wci_wci_cfwr_pw__whas ;
  assign WILL_FIRE_RL_wci_cfwr =
	     CAN_FIRE_RL_wci_cfwr && !WILL_FIRE_RL_wci_ctl_op_start &&
	     !WILL_FIRE_RL_wci_ctl_op_complete ;

  // rule RL_wci_ctlAckReg__dreg_update
  assign CAN_FIRE_RL_wci_ctlAckReg__dreg_update = 1'b1 ;
  assign WILL_FIRE_RL_wci_ctlAckReg__dreg_update = 1'b1 ;

  // rule RL_wci_respF_both
  assign CAN_FIRE_RL_wci_respF_both =
	     ((wci_respF_c_r == 2'b01) ?
		wci_respF_x_wire__whas :
		wci_respF_c_r != 2'b10 || wci_respF_x_wire__whas) &&
	     wci_respF_c_r != 2'b00 &&
	     wci_respF_enqueueing__whas ;
  assign WILL_FIRE_RL_wci_respF_both = CAN_FIRE_RL_wci_respF_both ;

  // rule RL_wci_respF_decCtr
  assign CAN_FIRE_RL_wci_respF_decCtr =
	     wci_respF_c_r != 2'b00 && !wci_respF_enqueueing__whas ;
  assign WILL_FIRE_RL_wci_respF_decCtr = CAN_FIRE_RL_wci_respF_decCtr ;

  // rule RL_wci_respF_incCtr
  assign CAN_FIRE_RL_wci_respF_incCtr =
	     ((wci_respF_c_r == 2'b00) ?
		wci_respF_x_wire__whas :
		wci_respF_c_r != 2'b01 || wci_respF_x_wire__whas) &&
	     wci_respF_enqueueing__whas &&
	     !(wci_respF_c_r != 2'b00) ;
  assign WILL_FIRE_RL_wci_respF_incCtr = CAN_FIRE_RL_wci_respF_incCtr ;

  // rule RL_wci_reqF__updateLevelCounter
  assign CAN_FIRE_RL_wci_reqF__updateLevelCounter =
	     (wci_wciReq__wget[59:57] != 3'b000) != wci_reqF_r_deq__whas ;
  assign WILL_FIRE_RL_wci_reqF__updateLevelCounter =
	     CAN_FIRE_RL_wci_reqF__updateLevelCounter ;

  // rule RL_mesgWF_portB
  assign CAN_FIRE_RL_mesgWF_portB = 1'b1 ;
  assign WILL_FIRE_RL_mesgWF_portB = 1'b1 ;

  // rule RL_mesgWF_portA
  assign CAN_FIRE_RL_mesgWF_portA = 1'b1 ;
  assign WILL_FIRE_RL_mesgWF_portA = 1'b1 ;

  // rule RL_wmemi_respAdvance
  assign CAN_FIRE_RL_wmemi_respAdvance =
	     wmemi_respF__FULL_N && wmemi_operateD && wmemi_peerIsReady &&
	     wmemi_wmemiResponse__wget[130:129] != 2'b00 ;
  assign WILL_FIRE_RL_wmemi_respAdvance = CAN_FIRE_RL_wmemi_respAdvance ;

  // rule RL_wmemi_peerIsReady__dreg_update
  assign CAN_FIRE_RL_wmemi_peerIsReady__dreg_update = 1'b1 ;
  assign WILL_FIRE_RL_wmemi_peerIsReady__dreg_update = 1'b1 ;

  // rule RL_wmemi_operateD__dreg_update
  assign CAN_FIRE_RL_wmemi_operateD__dreg_update = 1'b1 ;
  assign WILL_FIRE_RL_wmemi_operateD__dreg_update = 1'b1 ;

  // rule RL_wmemi_dhF_deq
  assign CAN_FIRE_RL_wmemi_dhF_deq = wmemiM_SDataAccept ;
  assign WILL_FIRE_RL_wmemi_dhF_deq = wmemiM_SDataAccept ;

  // rule RL_wmemi_reqF_deq
  assign CAN_FIRE_RL_wmemi_reqF_deq = wmemiM_SCmdAccept ;
  assign WILL_FIRE_RL_wmemi_reqF_deq = wmemiM_SCmdAccept ;

  // rule RL_wmemi_dhF_both
  assign CAN_FIRE_RL_wmemi_dhF_both =
	     ((wmemi_dhF_c_r == 2'b01) ?
		CAN_FIRE_RL_delay_write_req :
		wmemi_dhF_c_r != 2'b10 || CAN_FIRE_RL_delay_write_req) &&
	     wmemi_dhF_dequeueing__whas &&
	     CAN_FIRE_RL_delay_write_req ;
  assign WILL_FIRE_RL_wmemi_dhF_both = CAN_FIRE_RL_wmemi_dhF_both ;

  // rule RL_wmemi_dhF_decCtr
  assign CAN_FIRE_RL_wmemi_dhF_decCtr =
	     wmemi_dhF_dequeueing__whas && !CAN_FIRE_RL_delay_write_req ;
  assign WILL_FIRE_RL_wmemi_dhF_decCtr = CAN_FIRE_RL_wmemi_dhF_decCtr ;

  // rule RL_wmemi_dhF_incCtr
  assign CAN_FIRE_RL_wmemi_dhF_incCtr =
	     ((wmemi_dhF_c_r == 2'b00) ?
		CAN_FIRE_RL_delay_write_req :
		wmemi_dhF_c_r != 2'b01 || CAN_FIRE_RL_delay_write_req) &&
	     CAN_FIRE_RL_delay_write_req &&
	     !wmemi_dhF_dequeueing__whas ;
  assign WILL_FIRE_RL_wmemi_dhF_incCtr = CAN_FIRE_RL_wmemi_dhF_incCtr ;

  // rule RL_wmemi_reqF_both
  assign CAN_FIRE_RL_wmemi_reqF_both =
	     ((wmemi_reqF_c_r == 2'b01) ?
		wmemi_reqF_enqueueing__whas :
		wmemi_reqF_c_r != 2'b10 || wmemi_reqF_enqueueing__whas) &&
	     wmemi_reqF_dequeueing__whas &&
	     wmemi_reqF_enqueueing__whas ;
  assign WILL_FIRE_RL_wmemi_reqF_both = CAN_FIRE_RL_wmemi_reqF_both ;

  // rule RL_wmemi_reqF_incCtr
  assign CAN_FIRE_RL_wmemi_reqF_incCtr =
	     ((wmemi_reqF_c_r == 2'b00) ?
		wmemi_reqF_enqueueing__whas :
		wmemi_reqF_c_r != 2'b01 || wmemi_reqF_enqueueing__whas) &&
	     wmemi_reqF_enqueueing__whas &&
	     !wmemi_reqF_dequeueing__whas ;
  assign WILL_FIRE_RL_wmemi_reqF_incCtr = CAN_FIRE_RL_wmemi_reqF_incCtr ;

  // rule RL_wmemi_reqF_decCtr
  assign CAN_FIRE_RL_wmemi_reqF_decCtr =
	     wmemi_reqF_dequeueing__whas && !wmemi_reqF_enqueueing__whas ;
  assign WILL_FIRE_RL_wmemi_reqF_decCtr = CAN_FIRE_RL_wmemi_reqF_decCtr ;

  // inputs to muxes for submodule ports
  assign MUX_wci_illegalEdge__write_1__SEL_1 =
	     WILL_FIRE_RL_wci_ctl_op_complete && wci_illegalEdge ;
  assign MUX_wci_illegalEdge__write_1__VAL_2 =
	     wci_reqF__D_OUT[36:34] != 3'b100 && wci_reqF__D_OUT[36:34] != 3'b101 &&
	     wci_reqF__D_OUT[36:34] != 3'b110 ;
  assign MUX_wci_respF_c_r__write_1__VAL_2 = wci_respF_c_r + 2'b01 ;
  assign MUX_wci_respF_c_r__write_1__VAL_1 = wci_respF_c_r - 2'b01 ;
  assign MUX_wci_respF_x_wire__wset_1__VAL_2 =
	     wci_illegalEdge ? 34'h3C0DE4202 : 34'h1C0DE4201 ;
  assign MUX_wci_illegalEdge__write_1__SEL_2 =
	     WILL_FIRE_RL_wci_ctl_op_start &&
	     (wci_reqF__D_OUT[36:34] == 3'b000 && wci_cState != 3'b000 ||
	      wci_reqF__D_OUT[36:34] == 3'b001 && wci_cState != 3'b001 &&
	      wci_cState != 3'b011 ||
	      wci_reqF__D_OUT[36:34] == 3'b010 && wci_cState != 3'b010 ||
	      wci_reqF__D_OUT[36:34] == 3'b011 && wci_cState != 3'b011 &&
	      wci_cState != 3'b010 &&
	      wci_cState != 3'b001 ||
	      wci_reqF__D_OUT[36:34] == 3'b100 ||
	      wci_reqF__D_OUT[36:34] == 3'b101 ||
	      wci_reqF__D_OUT[36:34] == 3'b110 ||
	      wci_reqF__D_OUT[36:34] == 3'b111) ;
  assign MUX_wci_respF_q_0__write_1__SEL_2 =
	     WILL_FIRE_RL_wci_respF_incCtr && wci_respF_c_r == 2'b00 ;
  assign MUX_wci_respF_q_1__write_1__SEL_2 =
	     WILL_FIRE_RL_wci_respF_incCtr && wci_respF_c_r == 2'b01 ;
  assign MUX_wsiM_reqFifo_c_r__write_1__VAL_1 = wsiM_reqFifo_c_r - 2'b01 ;
  assign MUX_wsiM_reqFifo_c_r__write_1__VAL_2 = wsiM_reqFifo_c_r + 2'b01 ;
  assign MUX_wsiM_reqFifo_q_0__write_1__SEL_2 =
	     WILL_FIRE_RL_wsiM_reqFifo_incCtr && wsiM_reqFifo_c_r == 2'b00 ;
  assign MUX_wsiM_reqFifo_q_1__write_1__SEL_2 =
	     WILL_FIRE_RL_wsiM_reqFifo_incCtr && wsiM_reqFifo_c_r == 2'b01 ;
  assign MUX_mesgLength__write_1__VAL_2 =
	     (wsiS_reqFifo__D_OUT[39:8] == 32'b00000000000000000000000000000000) ?
	       15'b100000000000000 :
	       { 1'b1, wsiS_reqFifo__D_OUT[304:296], 5'b00000 } ;
  assign MUX_mesgLengthSoFar__write_1__VAL_2 = mesgLengthSoFar + 14'b00000000000001 ;
  assign MUX_opcode__write_1__VAL_2 = { 1'b1, wsiS_reqFifo__D_OUT[7:0] } ;
  assign MUX_unrollCnt__write_1__VAL_1 =
	     (metaRF__D_OUT[23:0] == 24'b000000000000000000000000) ? 16'b0000000000000001 : metaRF__D_OUT[20:5] ;
  assign MUX_unrollCnt__write_1__VAL_2 = unrollCnt - 16'b0000000000000001 ;
  assign MUX_wsiWordsRemain__write_1__VAL_2 = wsiWordsRemain - 12'b01 ;
  assign MUX_mesgLength__write_1__VAL_3 = { 1'b1, mlp1__h17953[8:0], 5'b00000 } ;
  assign MUX_mesgRdCount__write_1__SEL_1 =
	     WILL_FIRE_RL_wmrd_mesgBodyResponse && unrollCnt == 16'b0000000000000001 ;
  assign MUX_dlyRAG__write_1__VAL_1 = dlyRAG + 20'b00000000000000000001 ;
  assign MUX_dlyWAG__write_1__VAL_1 = dlyWAG + 20'b00000000000000000001 ;
  assign MUX_mesgRdCount__write_1__VAL_1 = mesgRdCount + 32'b00000000000000000000000000000001 ;
  assign MUX_mesgWtCount__write_1__VAL_1 = mesgWtCount + 32'b00000000000000000000000000000001 ;
  assign MUX_metaWF__enq_1__VAL_1 = { x1_opcode__h17253, x1_length__h17254 } ;
  assign MUX_rdSerPos__write_1__VAL_1 = rdSerPos + 2'b01 ;
  assign MUX_rdSerUnroll__write_1__VAL_2 = rdSerUnroll - 16'b0000000000000001 ;
  assign MUX_rdSyncWord__write_1__VAL_1 =
	     rdSerPos != 2'b11 && rdSerUnroll == 16'b0000000000000001 ;
  assign MUX_wmemi_dhF_c_r__write_1__VAL_1 = wmemi_dhF_c_r - 2'b01 ;
  assign MUX_wmemi_dhF_c_r__write_1__VAL_2 = wmemi_dhF_c_r + 2'b01 ;
  assign MUX_wmemi_dhF_q_0__write_1__VAL_2 =
	     { 2'b11, wide16Fa__D_OUT, 16'b1111111111111111 } ;
  assign MUX_wmemi_dhF_q_0__write_1__VAL_1 =
	     (wmemi_dhF_c_r == 2'b01) ?
	       MUX_wmemi_dhF_q_0__write_1__VAL_2 :
	       wmemi_dhF_q_1 ;
  assign MUX_wmemi_dhF_q_1__write_1__VAL_1 =
	     (wmemi_dhF_c_r == 2'b10) ?
	       MUX_wmemi_dhF_q_0__write_1__VAL_2 :
	       146'h0AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA ;
  assign MUX_wmemi_reqF_c_r__write_1__VAL_1 = wmemi_reqF_c_r - 2'b01 ;
  assign MUX_wmemi_reqF_c_r__write_1__VAL_2 = wmemi_reqF_c_r + 2'b01 ;
  assign MUX_wrtSerUnroll__write_1__VAL_1 = wrtSerUnroll - 16'b0000000000000001 ;
  assign MUX_wmemi_dhF_q_0__write_1__SEL_2 =
	     WILL_FIRE_RL_wmemi_dhF_incCtr && wmemi_dhF_c_r == 2'b00 ;
  assign MUX_wmemi_dhF_q_1__write_1__SEL_2 =
	     WILL_FIRE_RL_wmemi_dhF_incCtr && wmemi_dhF_c_r == 2'b01 ;
  assign MUX_wmemi_reqF_x_wire__wset_1__VAL_1 = { 4'b0101, addr__h20994, 12'b01 } ;
  assign MUX_wmemi_reqF_x_wire__wset_1__VAL_2 = { 4'b0011, addr__h21166, 12'b01 } ;
  assign MUX_wci_respF_x_wire__wset_1__VAL_1 = { 2'b01, x_data__h21804 } ;
  always@(WILL_FIRE_RL_wci_cfrd or
	  MUX_wci_respF_x_wire__wset_1__VAL_1 or
	  WILL_FIRE_RL_wci_ctl_op_complete or
	  MUX_wci_respF_x_wire__wset_1__VAL_2 or WILL_FIRE_RL_wci_cfwr)
  begin
    case (1'b1) // synopsys parallel_case
      WILL_FIRE_RL_wci_cfrd:
	  MUX_wci_respF_q_0__write_1__VAL_2 =
	      MUX_wci_respF_x_wire__wset_1__VAL_1;
      WILL_FIRE_RL_wci_ctl_op_complete:
	  MUX_wci_respF_q_0__write_1__VAL_2 =
	      MUX_wci_respF_x_wire__wset_1__VAL_2;
      WILL_FIRE_RL_wci_cfwr: MUX_wci_respF_q_0__write_1__VAL_2 = 34'h1C0DE4201;
      default: MUX_wci_respF_q_0__write_1__VAL_2 =
		   34'h2AAAAAAAA /* unspecified value */ ;
    endcase
  end
  assign MUX_wci_respF_q_0__write_1__VAL_1 =
	     (wci_respF_c_r == 2'b01) ?
	       MUX_wci_respF_q_0__write_1__VAL_2 :
	       wci_respF_q_1 ;
  assign MUX_wci_respF_q_1__write_1__VAL_1 =
	     (wci_respF_c_r == 2'b10) ?
	       MUX_wci_respF_q_0__write_1__VAL_2 :
	       34'h0AAAAAAAA ;
  assign MUX_rdSyncWord__write_1__VAL_2 =
	     rdSerPos != 2'b11 && v__h22720[23:0] == 24'b000000000000000000000000 ;
  assign MUX_wsiM_reqFifo_x_wire__wset_1__VAL_1 =
	     { 3'b001,
	       unrollCnt == 16'b0000000000000001,
	       1'b1,
	       x_burstLength__h22437,
	       mesg__h22346,
	       x_byteEn__h22438,
	       readMeta[31:24] } ;
  assign MUX_wsiM_reqFifo_q_0__write_1__VAL_2 =
	     WILL_FIRE_RL_wmrd_mesgBodyResponse ?
	       MUX_wsiM_reqFifo_x_wire__wset_1__VAL_1 :
	       wsiS_reqFifo__D_OUT ;
  assign MUX_wsiM_reqFifo_q_0__write_1__VAL_1 =
	     (wsiM_reqFifo_c_r == 2'b01) ?
	       MUX_wsiM_reqFifo_q_0__write_1__VAL_2 :
	       wsiM_reqFifo_q_1 ;
  assign MUX_wsiM_reqFifo_q_1__write_1__VAL_1 =
	     (wsiM_reqFifo_c_r == 2'b10) ?
	       MUX_wsiM_reqFifo_q_0__write_1__VAL_2 :
	       313'h00000AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA00 ;
  assign MUX_rdSerEmpty__write_1__PSEL_1 =
	     WILL_FIRE_RL_rdSer_begin || WILL_FIRE_RL_rdSer_body ;
  assign MUX_rdSerEmpty__write_1__SEL_1 =
	     MUX_rdSerEmpty__write_1__PSEL_1 &&
	     (rdSerEmpty || rdSerPos == 2'b00) ;
  assign MUX_dlyReadCredit_value__write_1__VAL_2 =
	     dlyReadCredit_value +
	     (WILL_FIRE_RL_delay_read_req ? 8'b11111111 : 8'b00000000) +
	     (CAN_FIRE_RL_delay_read_resp ? 8'b00000001 : 8'b00000000) ;
  assign MUX_dlyWordsStored_value__write_1__VAL_2 =
	     dlyWordsStored_value +
	     (CAN_FIRE_RL_delay_write_req ? 20'b00000000000000000001 : 20'b00000000000000000000) +
	     (WILL_FIRE_RL_delay_read_req ? 20'b00000000000000000001: 20'b00000000000000000000) ;
  assign MUX_wmemi_reqF_q_0__write_1__VAL_2 =
	     WILL_FIRE_RL_delay_read_req ?
	       MUX_wmemi_reqF_x_wire__wset_1__VAL_1 :
	       MUX_wmemi_reqF_x_wire__wset_1__VAL_2 ;
  assign MUX_wmemi_reqF_q_0__write_1__VAL_1 =
	     (wmemi_reqF_c_r == 2'b01) ?
	       MUX_wmemi_reqF_q_0__write_1__VAL_2 :
	       wmemi_reqF_q_1 ;
  assign MUX_wmemi_reqF_q_1__write_1__VAL_1 =
	     (wmemi_reqF_c_r == 2'b10) ?
	       MUX_wmemi_reqF_q_0__write_1__VAL_2 :
	       52'h0AAAAAAAAAAAA ;
  assign MUX_wmemi_reqF_q_0__write_1__SEL_2 =
	     WILL_FIRE_RL_wmemi_reqF_incCtr && wmemi_reqF_c_r == 2'b00 ;
  assign MUX_wmemi_reqF_q_1__write_1__SEL_2 =
	     WILL_FIRE_RL_wmemi_reqF_incCtr && wmemi_reqF_c_r == 2'b01 ;
  always@(wrtSerPos or
	  IF_wrtSerPos_11_EQ_2_14_THEN_0x0_ELSE_mesgWF_w_ETC___d354 or
	  x1__h19969 or x1__h19978)
  begin
    case (wrtSerPos)
      2'b00: MUX_wide16Fa__enq_1__VAL_2 = x1__h19969;
      2'b01: MUX_wide16Fa__enq_1__VAL_2 = x1__h19978;
      default: MUX_wide16Fa__enq_1__VAL_2 =
		   IF_wrtSerPos_11_EQ_2_14_THEN_0x0_ELSE_mesgWF_w_ETC___d354;
    endcase
  end
  always@(wrtSerPos or
	  IF_wrtSerPos_11_EQ_2_14_THEN_0x0_ELSE_metaWF_f_ETC___d377 or
	  x1__h20492 or x1__h20501)
  begin
    case (wrtSerPos)
      2'b00: MUX_wide16Fa__enq_1__VAL_1 = x1__h20492;
      2'b01: MUX_wide16Fa__enq_1__VAL_1 = x1__h20501;
      default: MUX_wide16Fa__enq_1__VAL_1 =
		   IF_wrtSerPos_11_EQ_2_14_THEN_0x0_ELSE_metaWF_f_ETC___d377;
    endcase
  end
  assign MUX_wrtSerPos__write_1__VAL_1 =
	     (wrtSerUnroll == 16'b0000000000000001) ? 2'b00 : wrtSerPos_11_PLUS_1___d1014 ;
  assign MUX_wrtSerPos__write_1__VAL_2 =
	     (metaWF__D_OUT[23:0] == 24'b000000000000000000000000) ?
	       2'b00 :
	       wrtSerPos_11_PLUS_1___d1014 ;
  assign MUX_endOfMessage__write_1__SEL_1 =
	     WILL_FIRE_RL_wmwt_messagePushImprecise &&
	     wsiS_reqFifo__D_OUT[307:296] == 12'b01 ;
  assign MUX_impreciseBurst__write_1__SEL_2 =
	     WILL_FIRE_RL_wmwt_mesgBegin && !wsiS_reqFifo__D_OUT[308] ;
  assign MUX_mesgLength__write_1__SEL_2 =
	     WILL_FIRE_RL_wmwt_mesgBegin && wsiS_reqFifo__D_OUT[308] ;
  assign MUX_metaWF__enq_1__SEL_1 =
	     WILL_FIRE_RL_wmwt_messageFinalize && impreciseBurst ;
  assign MUX_wrtSerStage__write_1__SEL_1 =
	     WILL_FIRE_RL_wrtSer_body && wrtSerPos == 2'b00 ;
  assign MUX_wrtSerStage_1__write_1__SEL_1 =
	     WILL_FIRE_RL_wrtSer_body && wrtSerPos == 2'b01 ;
  assign MUX_wrtSerStage_2__write_1__SEL_1 =
	     WILL_FIRE_RL_wrtSer_body && wrtSerPos == 2'b10 ;
  assign MUX_wrtSerStage_3__write_1__SEL_1 =
	     WILL_FIRE_RL_wrtSer_body && wrtSerPos == 2'b11 ;
  assign MUX_wide16Fa__enq_1__SEL_1 =
	     WILL_FIRE_RL_wrtSer_begin &&
	     (wrtSerPos == 2'b11 || metaWF__D_OUT[23:0] == 24'b000000000000000000000000) ;

  // inlined wires
  assign wci_wciReq__whas = 1'b1 ;
  assign wci_wciReq__wget =
	     { wciS0_MCmd,
	       wciS0_MAddrSpace,
	       wciS0_MByteEn,
	       wciS0_MAddr,
	       wciS0_MData } ;
  assign wci_reqF_r_enq__whas = CAN_FIRE_RL_wci_reqF_enq ;
  assign wci_reqF_r_clr__whas = 1'b0 ;
  assign wci_respF_dequeueing__whas = wci_respF_c_r != 2'b00 ;
  assign wci_wEdge__wget = wci_reqF__D_OUT[36:34] ;
  assign wci_sThreadBusy_pw__whas = 1'b0 ;
  assign wci_sFlagReg_1__wget = 1'b0 ;
  assign wci_wci_cfwr_pw__whas =
	     wci_reqF__EMPTY_N && wci_reqF__D_OUT[56] &&
	     wci_reqF__D_OUT[59:57] == 3'b001 ;
  assign wci_sFlagReg_1__whas = 1'b0 ;
  assign wci_wci_cfrd_pw__whas =
	     wci_reqF__EMPTY_N && wci_reqF__D_OUT[56] &&
	     wci_reqF__D_OUT[59:57] == 3'b010 ;
  assign wci_wci_ctrl_pw__whas =
	     wci_reqF__EMPTY_N && !wci_reqF__D_OUT[56] &&
	     wci_reqF__D_OUT[59:57] == 3'b010 ;
  assign wci_reqF_r_deq__whas =
	     WILL_FIRE_RL_wci_cfrd || WILL_FIRE_RL_wci_cfwr ||
	     WILL_FIRE_RL_wci_ctl_op_start ;
  assign wci_respF_enqueueing__whas =
	     WILL_FIRE_RL_wci_cfrd || WILL_FIRE_RL_wci_cfwr ||
	     WILL_FIRE_RL_wci_ctl_op_complete ;
  assign wci_respF_x_wire__whas =
	     WILL_FIRE_RL_wci_cfrd || WILL_FIRE_RL_wci_ctl_op_complete ||
	     WILL_FIRE_RL_wci_cfwr ;
  assign wci_wEdge__whas = WILL_FIRE_RL_wci_ctl_op_start ;
  assign wci_ctlAckReg_1__wget = 1'b1 ;
  assign wci_ctlAckReg_1__whas =
	     WILL_FIRE_RL_wci_ctrl_OrE || WILL_FIRE_RL_wci_ctrl_IsO ||
	     WILL_FIRE_RL_wci_ctrl_EiI ;
  assign wmemi_operateD_1__wget = 1'b1 ;
  assign wmemi_operateD_1__whas = wci_cState == 3'b010 ;
  assign wmemi_peerIsReady_1__whas = 1'b0 ;
  assign wmemi_peerIsReady_1__wget = 1'b0 ;
  assign wsiM_reqFifo_dequeueing__whas = CAN_FIRE_RL_wsiM_reqFifo_deq ;
  assign wsiM_sThreadBusy_pw__whas = wsiM1_SThreadBusy ;
  assign wsiM_operateD_1__wget = 1'b1 ;
  assign wsiM_operateD_1__whas = wci_cState == 3'b010 ;
  assign wsiM_peerIsReady_1__wget = 1'b1 ;
  assign wsiM_peerIsReady_1__whas = wsiM1_SReset_n ;
  assign wsiM_extStatusW__wget =
	     { wsiM_pMesgCount, wsiM_iMesgCount, wsiM_tBusyCount } ;
  assign wsiS_reqFifo_r_clr__whas = 1'b0 ;
  assign wsiS_wsiReq__wget =
	     { wsiS1_MCmd,
	       wsiS1_MReqLast,
	       wsiS1_MBurstPrecise,
	       wsiS1_MBurstLength,
	       wsiS1_MData,
	       wsiS1_MByteEn,
	       wsiS1_MReqInfo } ;
  assign wsiS_wsiReq__whas = 1'b1 ;
  assign wsiS_reqFifo_r_enq__whas = CAN_FIRE_RL_wsiS_reqFifo_enq ;
  assign wsiS_operateD_1__wget = 1'b1 ;
  assign wsiS_operateD_1__whas = wci_cState == 3'b010 ;
  assign wsiS_peerIsReady_1__wget = 1'b1 ;
  assign wsiS_peerIsReady_1__whas = wsiS1_MReset_n ;
  assign wsiS_extStatusW__wget =
	     { wsiS_pMesgCount, wsiS_iMesgCount, wsiS_tBusyCount } ;
  assign wsi_Es_mCmd_w__wget = wsiS1_MCmd ;
  assign wsi_Es_mCmd_w__whas = 1'b1 ;
  assign wsi_Es_mReqLast_w__whas = wsiS1_MReqLast ;
  assign wsi_Es_mBurstPrecise_w__whas = wsiS1_MBurstPrecise ;
  assign wsi_Es_mBurstLength_w__wget = wsiS1_MBurstLength ;
  assign wsi_Es_mBurstLength_w__whas = 1'b1 ;
  assign wsi_Es_mData_w__wget = wsiS1_MData ;
  assign wsi_Es_mData_w__whas = 1'b1 ;
  assign wsi_Es_mByteEn_w__whas = 1'b1 ;
  assign wsi_Es_mByteEn_w__wget = wsiS1_MByteEn ;
  assign wsi_Es_mReqInfo_w__wget = wsiS1_MReqInfo ;
  assign wsi_Es_mReqInfo_w__whas = 1'b1 ;
  assign wsi_Es_mDataInfo_w__whas = 1'b1 ;
  assign wsiM_reqFifo_enqueueing__whas =
	     WILL_FIRE_RL_wsipass_doMessagePush ||
	     WILL_FIRE_RL_wmrd_mesgBodyResponse ;
  assign wsiM_reqFifo_x_wire__whas =
	     WILL_FIRE_RL_wmrd_mesgBodyResponse ||
	     WILL_FIRE_RL_wsipass_doMessagePush ;
  assign wci_Es_mCmd_w__wget = wciS0_MCmd ;
  assign wci_Es_mCmd_w__whas = 1'b1 ;
  assign wci_Es_mAddrSpace_w__wget = wciS0_MAddrSpace ;
  assign wci_Es_mAddrSpace_w__whas = 1'b1 ;
  assign wci_Es_mAddr_w__wget = wciS0_MAddr ;
  assign wci_Es_mAddr_w__whas = 1'b1 ;
  assign wci_Es_mData_w__wget = wciS0_MData ;
  assign wci_Es_mByteEn_w__wget = wciS0_MByteEn ;
  assign wci_Es_mData_w__whas = 1'b1 ;
  assign wci_Es_mByteEn_w__whas = 1'b1 ;
  assign wmemi_reqF_dequeueing__whas =
	     wmemiM_SCmdAccept && wmemi_reqF_c_r != 2'b00 ;
  assign wmemi_dhF_enqueueing__whas = CAN_FIRE_RL_delay_write_req ;
  assign wmemi_dhF_x_wire__wget = MUX_wmemi_dhF_q_0__write_1__VAL_2 ;
  assign wmemi_dhF_x_wire__whas = CAN_FIRE_RL_delay_write_req ;
  assign wmemi_dhF_dequeueing__whas =
	     wmemiM_SDataAccept && wmemi_dhF_c_r != 2'b00 ;
  assign wmemi_wmemiResponse__wget =
	     { wmemiM_SResp, wmemiM_SRespLast, wmemiM_SData } ;
  assign wmemi_wmemiResponse__whas = 1'b1 ;
  assign wmemi_sDataAccept_w__wget = 1'b1 ;
  assign wmemi_sCmdAccept_w__wget = 1'b1 ;
  assign wmemi_sCmdAccept_w__whas = wmemiM_SCmdAccept ;
  assign wmemi_sDataAccept_w__whas = wmemiM_SDataAccept ;
  assign mesgWF_wDataIn__wget = wsiS_reqFifo__D_OUT[295:40] ;
  assign mesgWF_wDataOut__wget =
	     (mesgWF_rCache[267] && mesgWF_rCache[266:256] == mesgWF_rRdPtr) ?
	       mesgWF_rCache[255:0] :
	       mesgWF_memory__DOB ;
  assign mesgRF_wDataIn__whas = CAN_FIRE_RL_rdSer_body ;
  assign mesgWF_wDataOut__whas = 1'b1 ;
  assign mesgRF_pwDequeue__whas = CAN_FIRE_RL_wmrd_mesgBodyResponse ;
  assign mesgRF_pwEnqueue__whas = CAN_FIRE_RL_rdSer_body ;
  assign mesgRF_wDataOut__wget =
	     (mesgRF_rCache[267] && mesgRF_rCache[266:256] == mesgRF_rRdPtr) ?
	       mesgRF_rCache[255:0] :
	       mesgRF_memory__DOB ;
  assign mesgRF_wDataOut__whas = 1'b1 ;
  assign dlyWordsStored_acc_v1__wget = 20'b00000000000000000001 ;
  assign dlyWordsStored_acc_v1__whas = CAN_FIRE_RL_delay_write_req ;
  assign dlyWordsStored_acc_v2__wget = 20'b00000000000000000001 ;
  assign dlyReadCredit_acc_v1__wget = 8'b11111111 ;
  assign dlyReadCredit_acc_v2__wget = 8'b00000001 ;
  assign dlyReadCredit_acc_v2__whas = CAN_FIRE_RL_delay_read_resp ;
  assign wmemi_Em_sResp_w__wget = wmemiM_SResp ;
  assign wmemi_Em_sRespLast_w__whas = wmemiM_SRespLast ;
  assign wmemi_Em_sResp_w__whas = 1'b1 ;
  assign wmemi_Em_sData_w__wget = wmemiM_SData ;
  assign wmemi_Em_sData_w__whas = 1'b1 ;
  assign wci_respF_x_wire__wget = MUX_wci_respF_q_0__write_1__VAL_2 ;
  assign mesgRF_wDataIn__wget = { 224'b000000000000000000000000, v__h22720 } ;
  assign wsiM_reqFifo_x_wire__wget = MUX_wsiM_reqFifo_q_0__write_1__VAL_2 ;
  assign wmemi_reqF_enqueueing__whas =
	     WILL_FIRE_RL_delay_read_req || WILL_FIRE_RL_delay_write_req ;
  assign wmemi_reqF_x_wire__wget = MUX_wmemi_reqF_q_0__write_1__VAL_2 ;
  assign wmemi_reqF_x_wire__whas = wmemi_reqF_enqueueing__whas ;
  assign dlyWordsStored_acc_v2__whas = WILL_FIRE_RL_delay_read_req ;
  assign dlyReadCredit_acc_v1__whas = WILL_FIRE_RL_delay_read_req ;
  assign wsiS_reqFifo_r_deq__whas =
	     WILL_FIRE_RL_wsipass_doMessagePush ||
	     WILL_FIRE_RL_wmwt_messagePushPrecise ||
	     WILL_FIRE_RL_wmwt_messagePushImprecise ;
  assign mesgWF_pwEnqueue__whas =
	     WILL_FIRE_RL_wmwt_messagePushPrecise ||
	     WILL_FIRE_RL_wmwt_messagePushImprecise ;
  assign mesgWF_wDataIn__whas = mesgWF_pwEnqueue__whas ;
  assign mesgWF_pwDequeue__whas = CAN_FIRE_RL_wrtSer_body ;

  // register abortCount
  assign abortCount__D_IN = abortCount + 32'b00000000000000000000000000000001 ;
  assign abortCount__EN = CAN_FIRE_RL_wmwt_doAbort ;

  // register blockDelayWrite
  assign blockDelayWrite__D_IN =
	     WILL_FIRE_RL_delay_write_req && wrtDutyCount == 3'b111 ;
  assign blockDelayWrite__EN =
	     WILL_FIRE_RL_delay_write_req ||
	     WILL_FIRE_RL_delay_write_unblock ;

  // register bytesRead
  assign bytesRead__D_IN = bytesRead + 32'b00000000000000000000000000100000 ;
  assign bytesRead__EN =
	     MUX_rdSerEmpty__write_1__PSEL_1 && bytesRead != 32'hFFFFFFFF ;

  // register bytesWritten
  assign bytesWritten__D_IN = bytesWritten + 32'b00000000000000000000000000100000 ;
  assign bytesWritten__EN =
	     _dor1bytesWritten__EN_write && bytesWritten != 32'hFFFFFFFF ;

  // register cyclesPassed
  assign cyclesPassed__D_IN = cyclesPassed + 32'b000000000000000000000000001000001 ;
  assign cyclesPassed__EN = wsiS_statusR[0] && cyclesPassed != 32'hFFFFFFFF ;

  // register dlyCtrl
  assign dlyCtrl__D_IN = wci_reqF__D_OUT[31:0] ;
  assign dlyCtrl__EN =
	     WILL_FIRE_RL_wci_cfwr && wci_reqF__D_OUT[51:32] == 20'h0 ;

  // register dlyHoldoffBytes
  assign dlyHoldoffBytes__D_IN = wci_reqF__D_OUT[31:0] ;
  assign dlyHoldoffBytes__EN =
	     WILL_FIRE_RL_wci_cfwr && wci_reqF__D_OUT[51:32] == 20'h00004 ;

  // register dlyHoldoffCycles
  assign dlyHoldoffCycles__D_IN = wci_reqF__D_OUT[31:0] ;
  assign dlyHoldoffCycles__EN =
	     WILL_FIRE_RL_wci_cfwr && wci_reqF__D_OUT[51:32] == 20'h00008 ;

  // register dlyRAG
  assign dlyRAG__D_IN =
	     WILL_FIRE_RL_delay_read_req ? MUX_dlyRAG__write_1__VAL_1 : 20'b00000000000000000000 ;
  assign dlyRAG__EN =
	     WILL_FIRE_RL_delay_read_req || WILL_FIRE_RL_wci_ctrl_IsO ;

  // register dlyReadCredit_value
  assign dlyReadCredit_value__EN = 1'b1 ;
  assign dlyReadCredit_value__D_IN =
	     WILL_FIRE_RL_wci_ctrl_IsO ?
	       8'b00000001 :
	       MUX_dlyReadCredit_value__write_1__VAL_2 ;

  // register dlyWAG
  assign dlyWAG__D_IN =
	     WILL_FIRE_RL_delay_write_req ?
	       MUX_dlyWAG__write_1__VAL_1 :
	       20'b00000000000000000000 ;
  assign dlyWAG__EN =
	     WILL_FIRE_RL_delay_write_req || WILL_FIRE_RL_wci_ctrl_IsO ;

  // register dlyWordsStored_value
  assign dlyWordsStored_value__EN = 1'b1 ;
  assign dlyWordsStored_value__D_IN =
	     WILL_FIRE_RL_wci_ctrl_IsO ?
	       20'b00000000000000000000 :
	       MUX_dlyWordsStored_value__write_1__VAL_2 ;

  // register doAbort
  assign doAbort__D_IN = 1'b0 ;
  assign doAbort__EN = CAN_FIRE_RL_wmwt_doAbort ;

  // register endOfMessage
  assign endOfMessage__D_IN = MUX_endOfMessage__write_1__SEL_1 ;
  assign endOfMessage__EN =
	     WILL_FIRE_RL_wmwt_messagePushImprecise &&
	     wsiS_reqFifo__D_OUT[307:296] == 12'b01 ||
	     WILL_FIRE_RL_wmwt_messageFinalize ;

  // register errCount - jluu: removed because never used
//  assign errCount__D_IN = errCount + 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001 ;
//  assign errCount__EN =
//	     WILL_FIRE_RL_wmwt_messagePushImprecise &&
//	     wsiS_reqFifo__D_OUT[295:40] != valExpect &&
//	     (wsiS_reqFifo__D_OUT[307:296] != 12'b01 ||
//	      wsiS_reqFifo__D_OUT[39:8] != 32'b00000000000000000000000000000000) ;

  // register impreciseBurst
  always@(WILL_FIRE_RL_wmwt_doAbort or
	  MUX_impreciseBurst__write_1__SEL_2 or
	  WILL_FIRE_RL_wmwt_messageFinalize)
  case (1'b1)
    WILL_FIRE_RL_wmwt_doAbort: impreciseBurst__D_IN = 1'b0;
    MUX_impreciseBurst__write_1__SEL_2: impreciseBurst__D_IN = 1'b1;
    WILL_FIRE_RL_wmwt_messageFinalize: impreciseBurst__D_IN = 1'b0;
    default: impreciseBurst__D_IN = 1'b0 /* unspecified value */ ;
  endcase
  assign impreciseBurst__EN =
	     WILL_FIRE_RL_wmwt_mesgBegin && !wsiS_reqFifo__D_OUT[308] ||
	     WILL_FIRE_RL_wmwt_messageFinalize ||
	     WILL_FIRE_RL_wmwt_doAbort ;

  // register mesgLength
  always@(WILL_FIRE_RL_wmwt_doAbort or
	  MUX_mesgLength__write_1__SEL_2 or
	  MUX_mesgLength__write_1__VAL_2 or
	  MUX_endOfMessage__write_1__SEL_1 or
	  MUX_mesgLength__write_1__VAL_3 or WILL_FIRE_RL_wmwt_messageFinalize)
  case (1'b1)
    WILL_FIRE_RL_wmwt_doAbort: mesgLength__D_IN = 15'b010101010101010;
    MUX_mesgLength__write_1__SEL_2:
	mesgLength__D_IN = MUX_mesgLength__write_1__VAL_2;
    MUX_endOfMessage__write_1__SEL_1:
	mesgLength__D_IN = MUX_mesgLength__write_1__VAL_3;
    WILL_FIRE_RL_wmwt_messageFinalize: mesgLength__D_IN = 15'b010101010101010;
    default: mesgLength__D_IN = 15'b010101010101010 /* unspecified value */ ;
  endcase
  assign mesgLength__EN =
	     WILL_FIRE_RL_wmwt_messagePushImprecise &&
	     wsiS_reqFifo__D_OUT[307:296] == 12'b01 ||
	     WILL_FIRE_RL_wmwt_mesgBegin && wsiS_reqFifo__D_OUT[308] ||
	     WILL_FIRE_RL_wmwt_messageFinalize ||
	     WILL_FIRE_RL_wmwt_doAbort ;

  // register mesgLengthSoFar
  assign mesgLengthSoFar__D_IN =
	     MUX_impreciseBurst__write_1__SEL_2 ?
	       14'b00000000000000 :
	       MUX_mesgLengthSoFar__write_1__VAL_2 ;
  assign mesgLengthSoFar__EN =
	     WILL_FIRE_RL_wmwt_mesgBegin && !wsiS_reqFifo__D_OUT[308] ||
	     WILL_FIRE_RL_wmwt_messagePushImprecise ;

  // register mesgRF_rCache
  assign mesgRF_rCache__EN = CAN_FIRE_RL_rdSer_body ;
  assign mesgRF_rCache__D_IN = { 1'b1, mesgRF_rWrPtr, x__h16160 } ;

  // register mesgRF_rRdPtr
  assign mesgRF_rRdPtr__D_IN = x__h16052 ;
  assign mesgRF_rRdPtr__EN = CAN_FIRE_RL_wmrd_mesgBodyResponse ;

  // register mesgRF_rWrPtr
  assign mesgRF_rWrPtr__D_IN = mesgRF_rWrPtr + 11'b1 ;
  assign mesgRF_rWrPtr__EN = CAN_FIRE_RL_rdSer_body ;

  // register mesgRdCount
  assign mesgRdCount__D_IN =
	     MUX_mesgRdCount__write_1__SEL_1 ?
	       MUX_mesgRdCount__write_1__VAL_1 :
	       32'b00000000000000000000000000000000 ;
  assign mesgRdCount__EN =
	     WILL_FIRE_RL_wmrd_mesgBodyResponse && unrollCnt == 16'b0000000000000001 ||
	     WILL_FIRE_RL_wci_ctrl_IsO ;

  // register mesgReqValid
  assign mesgReqValid__D_IN = !WILL_FIRE_RL_wmwt_messageFinalize ;
  assign mesgReqValid__EN =
	     WILL_FIRE_RL_wmwt_messageFinalize ||
	     WILL_FIRE_RL_wmwt_requestPrecise ;

  // register mesgWF_rCache
  assign mesgWF_rCache__D_IN = { 1'b1, mesgWF_rWrPtr, x__h15234 } ;
  assign mesgWF_rCache__EN = mesgWF_pwEnqueue__whas ;

  // register mesgWF_rRdPtr
  assign mesgWF_rRdPtr__D_IN = x__h15126 ;
  assign mesgWF_rRdPtr__EN = CAN_FIRE_RL_wrtSer_body ;

  // register mesgWF_rWrPtr
  assign mesgWF_rWrPtr__D_IN = mesgWF_rWrPtr + 11'b1 ;
  assign mesgWF_rWrPtr__EN = mesgWF_pwEnqueue__whas ;

  // register mesgWtCount
  assign mesgWtCount__D_IN =
	     WILL_FIRE_RL_wmwt_messageFinalize ?
	       MUX_mesgWtCount__write_1__VAL_1 :
	       32'b00000000000000000000000000000000 ;
  assign mesgWtCount__EN =
	     WILL_FIRE_RL_wmwt_messageFinalize || WILL_FIRE_RL_wci_ctrl_IsO ;

  // register opcode
  always@(WILL_FIRE_RL_wmwt_doAbort or
	  WILL_FIRE_RL_wmwt_mesgBegin or
	  MUX_opcode__write_1__VAL_2 or WILL_FIRE_RL_wmwt_messageFinalize)
  case (1'b1)
    WILL_FIRE_RL_wmwt_doAbort: opcode__D_IN = 9'b010101010;
    WILL_FIRE_RL_wmwt_mesgBegin: opcode__D_IN = MUX_opcode__write_1__VAL_2;
    WILL_FIRE_RL_wmwt_messageFinalize: opcode__D_IN = 9'b010101010;
    default: opcode__D_IN = 9'b010101010 /* unspecified value */ ;
  endcase
  assign opcode__EN =
	     WILL_FIRE_RL_wmwt_messageFinalize || WILL_FIRE_RL_wmwt_doAbort ||
	     WILL_FIRE_RL_wmwt_mesgBegin ;

  // register preciseBurst
  always@(WILL_FIRE_RL_wmwt_doAbort or
	  MUX_mesgLength__write_1__SEL_2 or WILL_FIRE_RL_wmwt_messageFinalize)
  case (1'b1)
    WILL_FIRE_RL_wmwt_doAbort: preciseBurst__D_IN = 1'b0;
    MUX_mesgLength__write_1__SEL_2: preciseBurst__D_IN = 1'b1;
    WILL_FIRE_RL_wmwt_messageFinalize: preciseBurst__D_IN = 1'b0;
    default: preciseBurst__D_IN = 1'b0 /* unspecified value */ ;
  endcase
  assign preciseBurst__EN =
	     WILL_FIRE_RL_wmwt_mesgBegin && wsiS_reqFifo__D_OUT[308] ||
	     WILL_FIRE_RL_wmwt_messageFinalize ||
	     WILL_FIRE_RL_wmwt_doAbort ;

  // register rdSerAddr
  assign rdSerAddr__D_IN = 32'h0 ;
  assign rdSerAddr__EN = 1'b0 ;

  // register rdSerEmpty
  assign rdSerEmpty__D_IN = !MUX_rdSerEmpty__write_1__SEL_1 ;
  assign rdSerEmpty__EN =
	     (WILL_FIRE_RL_rdSer_begin || WILL_FIRE_RL_rdSer_body) &&
	     (rdSerEmpty || rdSerPos == 2'b00) ||
	     WILL_FIRE_RL_rdSer_sync ;

  // register rdSerMeta
  assign rdSerMeta__D_IN = metaRF__D_IN ;
  assign rdSerMeta__EN = CAN_FIRE_RL_rdSer_begin ;

  // register rdSerPos
  assign rdSerPos__D_IN =
	     MUX_rdSerEmpty__write_1__PSEL_1 ?
	       MUX_rdSerPos__write_1__VAL_1 :
	       2'b00 ;
  assign rdSerPos__EN =
	     WILL_FIRE_RL_rdSer_begin || WILL_FIRE_RL_rdSer_body ||
	     WILL_FIRE_RL_rdSer_sync ;

  // register rdSerStage
  assign rdSerStage__D_IN = wide16Fb__D_OUT[31:0] ;
  assign rdSerStage__EN =
	     MUX_rdSerEmpty__write_1__PSEL_1 &&
	     (rdSerEmpty || rdSerPos == 2'b00) ;

  // register rdSerStage_1
  assign rdSerStage_1__D_IN = wide16Fb__D_OUT[63:32] ;
  assign rdSerStage_1__EN =
	     MUX_rdSerEmpty__write_1__PSEL_1 &&
	     (rdSerEmpty || rdSerPos == 2'b00) ;

  // register rdSerStage_2
  assign rdSerStage_2__D_IN = wide16Fb__D_OUT[95:64] ;
  assign rdSerStage_2__EN =
	     MUX_rdSerEmpty__write_1__PSEL_1 &&
	     (rdSerEmpty || rdSerPos == 2'b00) ;

  // register rdSerStage_3
  assign rdSerStage_3__D_IN = wide16Fb__D_OUT[127:96] ;
  assign rdSerStage_3__EN =
	     MUX_rdSerEmpty__write_1__PSEL_1 &&
	     (rdSerEmpty || rdSerPos == 2'b00) ;

  // register rdSerUnroll
  assign rdSerUnroll__D_IN =
	     WILL_FIRE_RL_rdSer_begin ?
	       v__h22720[20:5] :
	       MUX_rdSerUnroll__write_1__VAL_2 ;
  assign rdSerUnroll__EN = MUX_rdSerEmpty__write_1__PSEL_1 ;

  // register rdSyncWord
  always@(WILL_FIRE_RL_rdSer_body or
	  MUX_rdSyncWord__write_1__VAL_1 or
	  WILL_FIRE_RL_rdSer_begin or
	  MUX_rdSyncWord__write_1__VAL_2 or WILL_FIRE_RL_rdSer_sync)
  begin
    case (1'b1) // synopsys parallel_case
      WILL_FIRE_RL_rdSer_body:
	  rdSyncWord__D_IN = MUX_rdSyncWord__write_1__VAL_1;
      WILL_FIRE_RL_rdSer_begin:
	  rdSyncWord__D_IN = MUX_rdSyncWord__write_1__VAL_2;
      WILL_FIRE_RL_rdSer_sync: rdSyncWord__D_IN = 1'b0;
      default: rdSyncWord__D_IN = 1'b0 /* unspecified value */ ;
    endcase
  end
  assign rdSyncWord__EN =
	     WILL_FIRE_RL_rdSer_body || WILL_FIRE_RL_rdSer_begin ||
	     WILL_FIRE_RL_rdSer_sync ;

  // register readMeta
  assign readMeta__D_IN = metaRF__D_OUT ;
  assign readMeta__EN = CAN_FIRE_RL_wmrd_mesgBegin ;

  // register readyToPush
  always@(WILL_FIRE_RL_wmwt_doAbort or
	  MUX_impreciseBurst__write_1__SEL_2 or
	  MUX_endOfMessage__write_1__SEL_1)
  case (1'b1)
    WILL_FIRE_RL_wmwt_doAbort: readyToPush__D_IN = 1'b0;
    MUX_impreciseBurst__write_1__SEL_2: readyToPush__D_IN = 1'b1;
    MUX_endOfMessage__write_1__SEL_1: readyToPush__D_IN = 1'b0;
    default: readyToPush__D_IN = 1'b0 /* unspecified value */ ;
  endcase
  assign readyToPush__EN =
	     WILL_FIRE_RL_wmwt_messagePushImprecise &&
	     wsiS_reqFifo__D_OUT[307:296] == 12'b01 ||
	     WILL_FIRE_RL_wmwt_mesgBegin && !wsiS_reqFifo__D_OUT[308] ||
	     WILL_FIRE_RL_wmwt_doAbort ;

  // register readyToRequest
  assign readyToRequest__D_IN = MUX_mesgLength__write_1__SEL_2 ;
  assign readyToRequest__EN =
	     WILL_FIRE_RL_wmwt_mesgBegin && wsiS_reqFifo__D_OUT[308] ||
	     WILL_FIRE_RL_wmwt_requestPrecise ;

  // register unrollCnt
  assign unrollCnt__D_IN =
	     WILL_FIRE_RL_wmrd_mesgBegin ?
	       MUX_unrollCnt__write_1__VAL_1 :
	       MUX_unrollCnt__write_1__VAL_2 ;
  assign unrollCnt__EN =
	     WILL_FIRE_RL_wmrd_mesgBegin ||
	     WILL_FIRE_RL_wmrd_mesgBodyResponse ;

  // register valExpect : jluu removed because never used
//  assign valExpect__D_IN = valExpect + 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001 ;
//  assign valExpect__EN =
//	     WILL_FIRE_RL_wmwt_messagePushImprecise &&
//	     (wsiS_reqFifo__D_OUT[307:296] != 12'b01 ||
//	      wsiS_reqFifo__D_OUT[39:8] != 32'b00000000000000000000000000000000) ;

  // register wci_cEdge
  assign wci_cEdge__D_IN = wci_reqF__D_OUT[36:34] ;
  assign wci_cEdge__EN = WILL_FIRE_RL_wci_ctl_op_start ;

  // register wci_cState
  assign wci_cState__D_IN = wci_nState ;
  assign wci_cState__EN =
	     WILL_FIRE_RL_wci_ctl_op_complete && !wci_illegalEdge ;

  // register wci_ctlAckReg
  assign wci_ctlAckReg__D_IN = wci_ctlAckReg_1__whas ;
  assign wci_ctlAckReg__EN = 1'b1 ;

  // register wci_ctlOpActive
  assign wci_ctlOpActive__D_IN = !WILL_FIRE_RL_wci_ctl_op_complete ;
  assign wci_ctlOpActive__EN =
	     WILL_FIRE_RL_wci_ctl_op_complete ||
	     WILL_FIRE_RL_wci_ctl_op_start ;

  // register wci_illegalEdge
  assign wci_illegalEdge__D_IN =
	     !MUX_wci_illegalEdge__write_1__SEL_1 &&
	     MUX_wci_illegalEdge__write_1__VAL_2 ;
  assign wci_illegalEdge__EN =
	     WILL_FIRE_RL_wci_ctl_op_complete && wci_illegalEdge ||
	     MUX_wci_illegalEdge__write_1__SEL_2 ;

  // register wci_nState
  always@(wci_reqF__D_OUT)
  begin
    case (wci_reqF__D_OUT[36:34])
      3'b000: wci_nState__D_IN = 3'b001;
      3'b001: wci_nState__D_IN = 3'b010;
      3'b010: wci_nState__D_IN = 3'b011;
      default: wci_nState__D_IN = 3'b000;
    endcase
  end
  assign wci_nState__EN =
	     WILL_FIRE_RL_wci_ctl_op_start &&
	     (wci_reqF__D_OUT[36:34] == 3'b000 && wci_cState == 3'b000 ||
	      wci_reqF__D_OUT[36:34] == 3'b001 &&
	      (wci_cState == 3'b001 || wci_cState == 3'b011) ||
	      wci_reqF__D_OUT[36:34] == 3'b010 && wci_cState == 3'b010 ||
	      wci_reqF__D_OUT[36:34] == 3'b011 &&
	      (wci_cState == 3'b011 || wci_cState == 3'b010 ||
	       wci_cState == 3'b001)) ;

  // register wci_reqF_countReg
  assign wci_reqF_countReg__D_IN =
	     (wci_wciReq__wget[59:57] != 3'b000) ?
	       wci_reqF_countReg + 2'b01 :
	       wci_reqF_countReg - 2'b01 ;
  assign wci_reqF_countReg__EN = CAN_FIRE_RL_wci_reqF__updateLevelCounter ;

  // register wci_respF_c_r
  assign wci_respF_c_r__D_IN =
	     WILL_FIRE_RL_wci_respF_decCtr ?
	       MUX_wci_respF_c_r__write_1__VAL_1 :
	       MUX_wci_respF_c_r__write_1__VAL_2 ;
  assign wci_respF_c_r__EN =
	     WILL_FIRE_RL_wci_respF_decCtr || WILL_FIRE_RL_wci_respF_incCtr ;

  // register wci_respF_q_0
  assign wci_respF_q_0__EN =
	     WILL_FIRE_RL_wci_respF_both ||
	     WILL_FIRE_RL_wci_respF_incCtr && wci_respF_c_r == 2'b00 ||
	     WILL_FIRE_RL_wci_respF_decCtr ;
  always@(WILL_FIRE_RL_wci_respF_both or
	  MUX_wci_respF_q_0__write_1__VAL_1 or
	  MUX_wci_respF_q_0__write_1__SEL_2 or
	  MUX_wci_respF_q_0__write_1__VAL_2 or
	  WILL_FIRE_RL_wci_respF_decCtr or wci_respF_q_1)
  begin
    case (1'b1) // synopsys parallel_case
      WILL_FIRE_RL_wci_respF_both:
	  wci_respF_q_0__D_IN = MUX_wci_respF_q_0__write_1__VAL_1;
      MUX_wci_respF_q_0__write_1__SEL_2:
	  wci_respF_q_0__D_IN = MUX_wci_respF_q_0__write_1__VAL_2;
      WILL_FIRE_RL_wci_respF_decCtr: wci_respF_q_0__D_IN = wci_respF_q_1;
      default: wci_respF_q_0__D_IN = 34'h2AAAAAAAA /* unspecified value */ ;
    endcase
  end

  // register wci_respF_q_1
  assign wci_respF_q_1__EN =
	     WILL_FIRE_RL_wci_respF_both ||
	     WILL_FIRE_RL_wci_respF_incCtr && wci_respF_c_r == 2'b01 ||
	     WILL_FIRE_RL_wci_respF_decCtr ;
  always@(WILL_FIRE_RL_wci_respF_both or
	  MUX_wci_respF_q_1__write_1__VAL_1 or
	  MUX_wci_respF_q_1__write_1__SEL_2 or
	  MUX_wci_respF_q_0__write_1__VAL_2 or WILL_FIRE_RL_wci_respF_decCtr)
  begin
    case (1'b1) // synopsys parallel_case
      WILL_FIRE_RL_wci_respF_both:
	  wci_respF_q_1__D_IN = MUX_wci_respF_q_1__write_1__VAL_1;
      MUX_wci_respF_q_1__write_1__SEL_2:
	  wci_respF_q_1__D_IN = MUX_wci_respF_q_0__write_1__VAL_2;
      WILL_FIRE_RL_wci_respF_decCtr: wci_respF_q_1__D_IN = 34'h0AAAAAAAA;
      default: wci_respF_q_1__D_IN = 34'h2AAAAAAAA /* unspecified value */ ;
    endcase
  end

  // register wci_sFlagReg
  assign wci_sFlagReg__D_IN = 1'b0 ;
  assign wci_sFlagReg__EN = 1'b1 ;

  // register wci_sThreadBusy_d
  assign wci_sThreadBusy_d__D_IN = 1'b0 ;
  assign wci_sThreadBusy_d__EN = 1'b1 ;

  // register wmemiRdReq
  assign wmemiRdReq__D_IN = wmemiRdReq + 32'b00000000000000000000000000000001 ;
  assign wmemiRdReq__EN = WILL_FIRE_RL_delay_read_req ;

  // register wmemiRdResp
  assign wmemiRdResp__D_IN = wmemiRdResp + 32'b00000000000000000000000000000001 ;
  assign wmemiRdResp__EN = CAN_FIRE_RL_delay_read_resp ;

  // register wmemiWrReq
  assign wmemiWrReq__D_IN = wmemiWrReq + 32'b00000000000000000000000000000001 ;
  assign wmemiWrReq__EN = CAN_FIRE_RL_delay_write_req ;

  // register wmemi_busyWithMessage
  assign wmemi_busyWithMessage__D_IN = 1'b0 ;
  assign wmemi_busyWithMessage__EN = 1'b0 ;

  // register wmemi_dhF_c_r
  assign wmemi_dhF_c_r__D_IN =
	     WILL_FIRE_RL_wmemi_dhF_decCtr ?
	       MUX_wmemi_dhF_c_r__write_1__VAL_1 :
	       MUX_wmemi_dhF_c_r__write_1__VAL_2 ;
  assign wmemi_dhF_c_r__EN =
	     WILL_FIRE_RL_wmemi_dhF_decCtr || WILL_FIRE_RL_wmemi_dhF_incCtr ;

  // register wmemi_dhF_q_0
  always@(WILL_FIRE_RL_wmemi_dhF_both or
	  MUX_wmemi_dhF_q_0__write_1__VAL_1 or
	  MUX_wmemi_dhF_q_0__write_1__SEL_2 or
	  MUX_wmemi_dhF_q_0__write_1__VAL_2 or
	  WILL_FIRE_RL_wmemi_dhF_decCtr or wmemi_dhF_q_1)
  begin
    case (1'b1) // synopsys parallel_case
      WILL_FIRE_RL_wmemi_dhF_both:
	  wmemi_dhF_q_0__D_IN = MUX_wmemi_dhF_q_0__write_1__VAL_1;
      MUX_wmemi_dhF_q_0__write_1__SEL_2:
	  wmemi_dhF_q_0__D_IN = MUX_wmemi_dhF_q_0__write_1__VAL_2;
      WILL_FIRE_RL_wmemi_dhF_decCtr: wmemi_dhF_q_0__D_IN = wmemi_dhF_q_1;
      default: wmemi_dhF_q_0__D_IN =
		   146'h2AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA /* unspecified value */ ;
    endcase
  end
  assign wmemi_dhF_q_0__EN =
	     WILL_FIRE_RL_wmemi_dhF_both ||
	     WILL_FIRE_RL_wmemi_dhF_incCtr && wmemi_dhF_c_r == 2'b00 ||
	     WILL_FIRE_RL_wmemi_dhF_decCtr ;

  // register wmemi_dhF_q_1
  always@(WILL_FIRE_RL_wmemi_dhF_both or
	  MUX_wmemi_dhF_q_1__write_1__VAL_1 or
	  MUX_wmemi_dhF_q_1__write_1__SEL_2 or
	  MUX_wmemi_dhF_q_0__write_1__VAL_2 or WILL_FIRE_RL_wmemi_dhF_decCtr)
  begin
    case (1'b1) // synopsys parallel_case
      WILL_FIRE_RL_wmemi_dhF_both:
	  wmemi_dhF_q_1__D_IN = MUX_wmemi_dhF_q_1__write_1__VAL_1;
      MUX_wmemi_dhF_q_1__write_1__SEL_2:
	  wmemi_dhF_q_1__D_IN = MUX_wmemi_dhF_q_0__write_1__VAL_2;
      WILL_FIRE_RL_wmemi_dhF_decCtr:
	  wmemi_dhF_q_1__D_IN = 146'h0AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
      default: wmemi_dhF_q_1__D_IN =
		   146'h2AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA /* unspecified value */ ;
    endcase
  end
  assign wmemi_dhF_q_1__EN =
	     WILL_FIRE_RL_wmemi_dhF_both ||
	     WILL_FIRE_RL_wmemi_dhF_incCtr && wmemi_dhF_c_r == 2'b01 ||
	     WILL_FIRE_RL_wmemi_dhF_decCtr ;

  // register wmemi_errorSticky
  assign wmemi_errorSticky__D_IN = 1'b0 ;
  assign wmemi_errorSticky__EN = 1'b0 ;

  // register wmemi_operateD
  assign wmemi_operateD__D_IN = wci_cState == 3'b010 ;
  assign wmemi_operateD__EN = 1'b1 ;

  // register wmemi_peerIsReady
  assign wmemi_peerIsReady__D_IN = 1'b1 ;
  assign wmemi_peerIsReady__EN = 1'b1 ;

  // register wmemi_reqF_c_r
  assign wmemi_reqF_c_r__D_IN =
	     WILL_FIRE_RL_wmemi_reqF_decCtr ?
	       MUX_wmemi_reqF_c_r__write_1__VAL_1 :
	       MUX_wmemi_reqF_c_r__write_1__VAL_2 ;
  assign wmemi_reqF_c_r__EN =
	     WILL_FIRE_RL_wmemi_reqF_decCtr ||
	     WILL_FIRE_RL_wmemi_reqF_incCtr ;

  // register wmemi_reqF_q_0
  always@(WILL_FIRE_RL_wmemi_reqF_both or
	  MUX_wmemi_reqF_q_0__write_1__VAL_1 or
	  MUX_wmemi_reqF_q_0__write_1__SEL_2 or
	  MUX_wmemi_reqF_q_0__write_1__VAL_2 or
	  WILL_FIRE_RL_wmemi_reqF_decCtr or wmemi_reqF_q_1)
  begin
    case (1'b1) // synopsys parallel_case
      WILL_FIRE_RL_wmemi_reqF_both:
	  wmemi_reqF_q_0__D_IN = MUX_wmemi_reqF_q_0__write_1__VAL_1;
      MUX_wmemi_reqF_q_0__write_1__SEL_2:
	  wmemi_reqF_q_0__D_IN = MUX_wmemi_reqF_q_0__write_1__VAL_2;
      WILL_FIRE_RL_wmemi_reqF_decCtr: wmemi_reqF_q_0__D_IN = wmemi_reqF_q_1;
      default: wmemi_reqF_q_0__D_IN =
		   52'hAAAAAAAAAAAAA /* unspecified value */ ;
    endcase
  end
  assign wmemi_reqF_q_0__EN =
	     WILL_FIRE_RL_wmemi_reqF_both ||
	     WILL_FIRE_RL_wmemi_reqF_incCtr && wmemi_reqF_c_r == 2'b00 ||
	     WILL_FIRE_RL_wmemi_reqF_decCtr ;

  // register wmemi_reqF_q_1
  always@(WILL_FIRE_RL_wmemi_reqF_both or
	  MUX_wmemi_reqF_q_1__write_1__VAL_1 or
	  MUX_wmemi_reqF_q_1__write_1__SEL_2 or
	  MUX_wmemi_reqF_q_0__write_1__VAL_2 or WILL_FIRE_RL_wmemi_reqF_decCtr)
  begin
    case (1'b1) // synopsys parallel_case
      WILL_FIRE_RL_wmemi_reqF_both:
	  wmemi_reqF_q_1__D_IN = MUX_wmemi_reqF_q_1__write_1__VAL_1;
      MUX_wmemi_reqF_q_1__write_1__SEL_2:
	  wmemi_reqF_q_1__D_IN = MUX_wmemi_reqF_q_0__write_1__VAL_2;
      WILL_FIRE_RL_wmemi_reqF_decCtr: wmemi_reqF_q_1__D_IN = 52'h0AAAAAAAAAAAA;
      default: wmemi_reqF_q_1__D_IN =
		   52'hAAAAAAAAAAAAA /* unspecified value */ ;
    endcase
  end
  assign wmemi_reqF_q_1__EN =
	     WILL_FIRE_RL_wmemi_reqF_both ||
	     WILL_FIRE_RL_wmemi_reqF_incCtr && wmemi_reqF_c_r == 2'b01 ||
	     WILL_FIRE_RL_wmemi_reqF_decCtr ;

  // register wmemi_statusR
  assign wmemi_statusR__D_IN =
	     { wmemi_isReset__VAL,
	       !wmemi_peerIsReady,
	       !wmemi_operateD,
	       wmemi_errorSticky,
	       3'b000,
	       wmemi_trafficSticky } ;
  assign wmemi_statusR__EN = 1'b1 ;

  // register wmemi_trafficSticky
  assign wmemi_trafficSticky__D_IN = 1'b1 ;
  assign wmemi_trafficSticky__EN = wmemiM_SCmdAccept ;

  // register wrtDutyCount
  assign wrtDutyCount__D_IN = wrtDutyCount + 3'b001 ;
  assign wrtDutyCount__EN = CAN_FIRE_RL_delay_write_req ;

  // register wrtSerAddr
  assign wrtSerAddr__D_IN = 32'h0 ;
  assign wrtSerAddr__EN = 1'b0 ;

  // register wrtSerMeta
  assign wrtSerMeta__D_IN = metaWF__D_OUT ;
  assign wrtSerMeta__EN = CAN_FIRE_RL_wrtSer_begin ;

  // register wrtSerPos
  assign wrtSerPos__D_IN =
	     WILL_FIRE_RL_wrtSer_body ?
	       MUX_wrtSerPos__write_1__VAL_1 :
	       MUX_wrtSerPos__write_1__VAL_2 ;
  assign wrtSerPos__EN =
	     WILL_FIRE_RL_wrtSer_body || WILL_FIRE_RL_wrtSer_begin ;

  // register wrtSerStage
  assign wrtSerStage__D_IN =
	     MUX_wrtSerStage__write_1__SEL_1 ? x__h19905[31:0] : metaWF__D_OUT ;
  assign wrtSerStage__EN =
	     WILL_FIRE_RL_wrtSer_body && wrtSerPos == 2'b00 ||
	     WILL_FIRE_RL_wrtSer_begin && wrtSerPos == 2'b00 ;

  // register wrtSerStage_1
  assign wrtSerStage_1__D_IN =
	     MUX_wrtSerStage_1__write_1__SEL_1 ?
	       x__h19905[31:0] :
	       metaWF__D_OUT ;
  assign wrtSerStage_1__EN =
	     WILL_FIRE_RL_wrtSer_body && wrtSerPos == 2'b01 ||
	     WILL_FIRE_RL_wrtSer_begin && wrtSerPos == 2'b01 ;

  // register wrtSerStage_2
  assign wrtSerStage_2__D_IN =
	     MUX_wrtSerStage_2__write_1__SEL_1 ?
	       x__h19905[31:0] :
	       metaWF__D_OUT ;
  assign wrtSerStage_2__EN =
	     WILL_FIRE_RL_wrtSer_body && wrtSerPos == 2'b10 ||
	     WILL_FIRE_RL_wrtSer_begin && wrtSerPos == 2'b10 ;

  // register wrtSerStage_3
  assign wrtSerStage_3__D_IN =
	     MUX_wrtSerStage_3__write_1__SEL_1 ?
	       x__h19905[31:0] :
	       metaWF__D_OUT ;
  assign wrtSerStage_3__EN =
	     WILL_FIRE_RL_wrtSer_body && wrtSerPos == 2'b11 ||
	     WILL_FIRE_RL_wrtSer_begin && wrtSerPos == 2'b11 ;

  // register wrtSerUnroll
  assign wrtSerUnroll__D_IN =
	     WILL_FIRE_RL_wrtSer_body ?
	       MUX_wrtSerUnroll__write_1__VAL_1 :
	       metaWF__D_OUT[20:5] ;
  assign wrtSerUnroll__EN =
	     WILL_FIRE_RL_wrtSer_body || WILL_FIRE_RL_wrtSer_begin ;

  // register wsiM_burstKind
  assign wsiM_burstKind__D_IN =
	     (wsiM_burstKind == 2'b00) ?
	       (wsiM_reqFifo_q_0[308] ? 2'b01 : 2'b10) :
	       2'b00 ;
  assign wsiM_burstKind__EN =
	     WILL_FIRE_RL_wsiM_reqFifo_deq &&
	     wsiM_reqFifo_q_0[312:310] == 3'b001 &&
	     (wsiM_burstKind == 2'b00 ||
	      wsiM_burstKind == 2'b01 && wsiM_reqFifo_q_0[309] ||
	      wsiM_burstKind == 2'b10 && wsiM_reqFifo_q_0[307:296] == 12'b01) ;

  // register wsiM_errorSticky
  assign wsiM_errorSticky__D_IN = 1'b0 ;
  assign wsiM_errorSticky__EN = 1'b0 ;

  // register wsiM_iMesgCount
  assign wsiM_iMesgCount__D_IN = wsiM_iMesgCount + 32'b00000000000000000000000000000001 ;
  assign wsiM_iMesgCount__EN =
	     WILL_FIRE_RL_wsiM_reqFifo_deq &&
	     wsiM_reqFifo_q_0[312:310] == 3'b001 &&
	     wsiM_burstKind == 2'b10 &&
	     wsiM_reqFifo_q_0[307:296] == 12'b01 ;

  // register wsiM_operateD
  assign wsiM_operateD__D_IN = wci_cState == 3'b010 ;
  assign wsiM_operateD__EN = 1'b1 ;

  // register wsiM_pMesgCount
  assign wsiM_pMesgCount__D_IN = wsiM_pMesgCount + 32'b00000000000000000000000000000001;
  assign wsiM_pMesgCount__EN =
	     WILL_FIRE_RL_wsiM_reqFifo_deq &&
	     wsiM_reqFifo_q_0[312:310] == 3'b001 &&
	     wsiM_burstKind == 2'b01 &&
	     wsiM_reqFifo_q_0[309] ;

  // register wsiM_peerIsReady
  assign wsiM_peerIsReady__D_IN = wsiM1_SReset_n ;
  assign wsiM_peerIsReady__EN = 1'b1 ;

  // register wsiM_reqFifo_c_r
  assign wsiM_reqFifo_c_r__D_IN =
	     WILL_FIRE_RL_wsiM_reqFifo_decCtr ?
	       MUX_wsiM_reqFifo_c_r__write_1__VAL_1 :
	       MUX_wsiM_reqFifo_c_r__write_1__VAL_2 ;
  assign wsiM_reqFifo_c_r__EN =
	     WILL_FIRE_RL_wsiM_reqFifo_decCtr ||
	     WILL_FIRE_RL_wsiM_reqFifo_incCtr ;

  // register wsiM_reqFifo_q_0
  assign wsiM_reqFifo_q_0__EN =
	     WILL_FIRE_RL_wsiM_reqFifo_both ||
	     WILL_FIRE_RL_wsiM_reqFifo_incCtr && wsiM_reqFifo_c_r == 2'b00 ||
	     WILL_FIRE_RL_wsiM_reqFifo_decCtr ;
  always@(WILL_FIRE_RL_wsiM_reqFifo_both or
	  MUX_wsiM_reqFifo_q_0__write_1__VAL_1 or
	  MUX_wsiM_reqFifo_q_0__write_1__SEL_2 or
	  MUX_wsiM_reqFifo_q_0__write_1__VAL_2 or
	  WILL_FIRE_RL_wsiM_reqFifo_decCtr or wsiM_reqFifo_q_1)
  begin
    case (1'b1) // synopsys parallel_case
      WILL_FIRE_RL_wsiM_reqFifo_both:
	  wsiM_reqFifo_q_0__D_IN = MUX_wsiM_reqFifo_q_0__write_1__VAL_1;
      MUX_wsiM_reqFifo_q_0__write_1__SEL_2:
	  wsiM_reqFifo_q_0__D_IN = MUX_wsiM_reqFifo_q_0__write_1__VAL_2;
      WILL_FIRE_RL_wsiM_reqFifo_decCtr:
	  wsiM_reqFifo_q_0__D_IN = wsiM_reqFifo_q_1;
      default: wsiM_reqFifo_q_0__D_IN =
		   313'h0AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA /* unspecified value */ ;
    endcase
  end

  // register wsiM_reqFifo_q_1
  assign wsiM_reqFifo_q_1__EN =
	     WILL_FIRE_RL_wsiM_reqFifo_both ||
	     WILL_FIRE_RL_wsiM_reqFifo_incCtr && wsiM_reqFifo_c_r == 2'b01 ||
	     WILL_FIRE_RL_wsiM_reqFifo_decCtr ;
  always@(WILL_FIRE_RL_wsiM_reqFifo_both or
	  MUX_wsiM_reqFifo_q_1__write_1__VAL_1 or
	  MUX_wsiM_reqFifo_q_1__write_1__SEL_2 or
	  MUX_wsiM_reqFifo_q_0__write_1__VAL_2 or
	  WILL_FIRE_RL_wsiM_reqFifo_decCtr)
  begin
    case (1'b1) // synopsys parallel_case
      WILL_FIRE_RL_wsiM_reqFifo_both:
	  wsiM_reqFifo_q_1__D_IN = MUX_wsiM_reqFifo_q_1__write_1__VAL_1;
      MUX_wsiM_reqFifo_q_1__write_1__SEL_2:
	  wsiM_reqFifo_q_1__D_IN = MUX_wsiM_reqFifo_q_0__write_1__VAL_2;
      WILL_FIRE_RL_wsiM_reqFifo_decCtr:
	  wsiM_reqFifo_q_1__D_IN =
	      313'h00000AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA00;
      default: wsiM_reqFifo_q_1__D_IN =
		   313'h0AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA /* unspecified value */ ;
    endcase
  end

  // register wsiM_sThreadBusy_d
  assign wsiM_sThreadBusy_d__D_IN = wsiM1_SThreadBusy ;
  assign wsiM_sThreadBusy_d__EN = 1'b1 ;

  // register wsiM_statusR
  assign wsiM_statusR__D_IN =
	     { wsiM_isReset__VAL,
	       !wsiM_peerIsReady,
	       !wsiM_operateD,
	       wsiM_errorSticky,
	       wsiM_burstKind != 2'b00,
	       wsiM_sThreadBusy_d,
	       1'b0,
	       wsiM_trafficSticky } ;
  assign wsiM_statusR__EN = 1'b1 ;

  // register wsiM_tBusyCount
  assign wsiM_tBusyCount__D_IN = wsiM_tBusyCount + 32'b00000000000000000000000000000001 ;
  assign wsiM_tBusyCount__EN = CAN_FIRE_RL_wsiM_inc_tBusyCount ;

  // register wsiM_trafficSticky
  assign wsiM_trafficSticky__D_IN = 1'b1 ;
  assign wsiM_trafficSticky__EN =
	     WILL_FIRE_RL_wsiM_reqFifo_deq &&
	     wsiM_reqFifo_q_0[312:310] == 3'b001 ;

  // register wsiS_burstKind
  assign wsiS_burstKind__D_IN =
	     (wsiS_burstKind == 2'b00) ?
	       (wsiS_wsiReq__wget[308] ? 2'b01 : 2'b10) :
	       2'b00 ;
  assign wsiS_burstKind__EN =
	     WILL_FIRE_RL_wsiS_reqFifo_enq &&
	     (wsiS_burstKind == 2'b00 ||
	      wsiS_burstKind == 2'b01 && wsiS_wsiReq__wget[309] ||
	      wsiS_burstKind == 2'b10 && wsiS_wsiReq__wget[307:296] == 12'b01) ;

  // register wsiS_errorSticky
  assign wsiS_errorSticky__D_IN = 1'b1 ;
  assign wsiS_errorSticky__EN =
	     WILL_FIRE_RL_wsiS_reqFifo_enq && !wsiS_reqFifo__FULL_N ;

  // register wsiS_iMesgCount
  assign wsiS_iMesgCount__D_IN = wsiS_iMesgCount + 32'b00000000000000000000000000000001 ;
  assign wsiS_iMesgCount__EN =
	     WILL_FIRE_RL_wsiS_reqFifo_enq && wsiS_burstKind == 2'b10 &&
	     wsiS_wsiReq__wget[307:296] == 12'b01 ;

  // register wsiS_operateD
  assign wsiS_operateD__D_IN = wci_cState == 3'b010 ;
  assign wsiS_operateD__EN = 1'b1 ;

  // register wsiS_pMesgCount
  assign wsiS_pMesgCount__D_IN = wsiS_pMesgCount + 32'b00000000000000000000000000000001 ;
  assign wsiS_pMesgCount__EN =
	     WILL_FIRE_RL_wsiS_reqFifo_enq && wsiS_burstKind == 2'b01 &&
	     wsiS_wsiReq__wget[309] ;

  // register wsiS_peerIsReady
  assign wsiS_peerIsReady__D_IN = wsiS1_MReset_n ;
  assign wsiS_peerIsReady__EN = 1'b1 ;

  // register wsiS_reqFifo_countReg
  assign wsiS_reqFifo_countReg__D_IN =
	     CAN_FIRE_RL_wsiS_reqFifo_enq ?
	       wsiS_reqFifo_countReg + 2'b01 :
	       wsiS_reqFifo_countReg - 2'b01 ;
  assign wsiS_reqFifo_countReg__EN =
	     CAN_FIRE_RL_wsiS_reqFifo__updateLevelCounter ;

  // register wsiS_statusR
  assign wsiS_statusR__EN = 1'b1 ;
  assign wsiS_statusR__D_IN =
	     { wsiS_isReset__VAL,
	       !wsiS_peerIsReady,
	       !wsiS_operateD,
	       wsiS_errorSticky,
	       wsiS_burstKind != 2'b00,
	       NOT_wsiS_reqFifo_countReg_96_ULE_1_97___d698 ||
	       wsiS_isReset__VAL ||
	       !wsiS_operateD ||
	       !wsiS_peerIsReady,
	       1'b0,
	       wsiS_trafficSticky } ;

  // register wsiS_tBusyCount
  assign wsiS_tBusyCount__D_IN = wsiS_tBusyCount + 32'b00000000000000000000000000000001 ;
  assign wsiS_tBusyCount__EN = CAN_FIRE_RL_wsiS_inc_tBusyCount ;

  // register wsiS_trafficSticky
  assign wsiS_trafficSticky__D_IN = 1'b1 ;
  assign wsiS_trafficSticky__EN = CAN_FIRE_RL_wsiS_reqFifo_enq ;

  // register wsiWordsRemain
  assign wsiWordsRemain__D_IN =
	     MUX_mesgLength__write_1__SEL_2 ?
	       wsiS_reqFifo__D_OUT[307:296] :
	       MUX_wsiWordsRemain__write_1__VAL_2 ;
  assign wsiWordsRemain__EN =
	     WILL_FIRE_RL_wmwt_mesgBegin && wsiS_reqFifo__D_OUT[308] ||
	     WILL_FIRE_RL_wmwt_messagePushPrecise ;

  // register zeroLengthMesg
  assign zeroLengthMesg__D_IN = wsiS_reqFifo__D_OUT[39:8] == 32'b00000000000000000000000000000000 ;
  assign zeroLengthMesg__EN = MUX_mesgLength__write_1__SEL_2 ;

  // submodule mesgRF_memory
  assign mesgRF_memory__WEA = CAN_FIRE_RL_rdSer_body ;
  assign mesgRF_memory__ADDRA = mesgRF_rWrPtr[9:0] ;
  assign mesgRF_memory__WEB = 1'b0 ;
  assign mesgRF_memory__ADDRB =
	     CAN_FIRE_RL_wmrd_mesgBodyResponse ?
	       x__h16052[9:0] :
	       mesgRF_rRdPtr[9:0] ;
  assign mesgRF_memory__DIB =
	     256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA /* unspecified value */  ;
  assign mesgRF_memory__ENA = 1'b1 ;
  assign mesgRF_memory__ENB = 1'b1 ;
  assign mesgRF_memory__DIA = x__h16160 ;

  // submodule mesgWF_memory
  assign mesgWF_memory__ADDRA = mesgWF_rWrPtr[9:0] ;
  assign mesgWF_memory__WEB = 1'b0 ;
  assign mesgWF_memory__DIB =
	     256'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA /* unspecified value */  ;
  assign mesgWF_memory__ENA = 1'b1 ;
  assign mesgWF_memory__ENB = 1'b1 ;
  assign mesgWF_memory__WEA = mesgWF_pwEnqueue__whas ;
  assign mesgWF_memory__DIA = x__h15234 ;
  assign mesgWF_memory__ADDRB =
	     CAN_FIRE_RL_wrtSer_body ? x__h15126[9:0] : mesgWF_rRdPtr[9:0] ;

  // submodule metaRF
  always@(rdSerPos or
	  rdSerStage_3 or wide16Fb__D_OUT or rdSerStage_1 or rdSerStage_2)
  begin
    case (rdSerPos)
      2'b00: metaRF__D_IN = wide16Fb__D_OUT[31:0];
      2'b01: metaRF__D_IN = rdSerStage_1;
      2'b10: metaRF__D_IN = rdSerStage_2;
      2'b11: metaRF__D_IN = rdSerStage_3;
    endcase
  end
  assign metaRF__DEQ = CAN_FIRE_RL_wmrd_mesgBegin ;
  assign metaRF__CLR = 1'b0 ;
  assign metaRF__ENQ = CAN_FIRE_RL_rdSer_begin ;

  // submodule metaWF
  assign metaWF__CLR = 1'b0 ;
  assign metaWF__D_IN =
	     MUX_metaWF__enq_1__SEL_1 ?
	       MUX_metaWF__enq_1__VAL_1 :
	       MUX_metaWF__enq_1__VAL_1 ;
  assign metaWF__ENQ =
	     WILL_FIRE_RL_wmwt_messageFinalize && impreciseBurst ||
	     WILL_FIRE_RL_wmwt_requestPrecise ;
  assign metaWF__DEQ = CAN_FIRE_RL_wrtSer_begin ;

  // submodule wci_reqF
  assign wci_reqF__D_IN = wci_wciReq__wget ;
  assign wci_reqF__DEQ = wci_reqF_r_deq__whas ;
  assign wci_reqF__ENQ = CAN_FIRE_RL_wci_reqF_enq ;
  assign wci_reqF__CLR = 1'b0 ;

  // submodule wide16Fa
  assign wide16Fa__DEQ = CAN_FIRE_RL_delay_write_req ;
  assign wide16Fa__CLR = 1'b0 ;
  assign wide16Fa__D_IN =
	     MUX_wide16Fa__enq_1__SEL_1 ?
	       MUX_wide16Fa__enq_1__VAL_1 :
	       MUX_wide16Fa__enq_1__VAL_2 ;
  assign wide16Fa__ENQ =
	     WILL_FIRE_RL_wrtSer_begin &&
	     (wrtSerPos == 2'b11 || metaWF__D_OUT[23:0] == 24'b000000000000000000000000) ||
	     WILL_FIRE_RL_wrtSer_body &&
	     (wrtSerPos == 2'b11 || wrtSerUnroll == 16'b0000000000000001) ;

  // submodule wide16Fb
  assign wide16Fb__D_IN = wmemi_respF__D_OUT[127:0] ;
  assign wide16Fb__ENQ = CAN_FIRE_RL_delay_read_resp ;
  assign wide16Fb__CLR = 1'b0 ;
  assign wide16Fb__DEQ =
	     MUX_rdSerEmpty__write_1__PSEL_1 &&
	     (rdSerEmpty || rdSerPos == 2'b00) ;

  // submodule wmemi_respF
  assign wmemi_respF__D_IN = wmemi_wmemiResponse__wget ;
  assign wmemi_respF__DEQ = CAN_FIRE_RL_delay_read_resp ;
  assign wmemi_respF__ENQ = CAN_FIRE_RL_wmemi_respAdvance ;
  assign wmemi_respF__CLR = 1'b0 ;

  // submodule wsiS_reqFifo
  assign wsiS_reqFifo__D_IN = wsiS_wsiReq__wget ;
  assign wsiS_reqFifo__ENQ = CAN_FIRE_RL_wsiS_reqFifo_enq ;
  assign wsiS_reqFifo__CLR = 1'b0 ;
  assign wsiS_reqFifo__DEQ = wsiS_reqFifo_r_deq__whas ;

  // remaining internal signals
  assign IF_wrtSerPos_11_EQ_2_14_THEN_0x0_ELSE_mesgWF_w_ETC___d354 =
	     { (wrtSerPos == 2'b10) ? 32'h0 : x__h19905[31:0],
	       (wrtSerPos == 2'b10) ? x__h19905[31:0] : wrtSerStage_2,
	       wrtSerStage_1,
	       wrtSerStage } ;
  assign IF_wrtSerPos_11_EQ_2_14_THEN_0x0_ELSE_metaWF_f_ETC___d377 =
	     { (wrtSerPos == 2'b10) ? 32'h0 : metaWF__D_OUT,
	       (wrtSerPos == 2'b10) ? metaWF__D_OUT : wrtSerStage_2,
	       wrtSerStage_1,
	       wrtSerStage } ;
  assign NOT_dlyWordsStored_value_13_SLE_0_64_65_AND_NO_ETC___d272 =
	     (dlyWordsStored_value ^ 20'h80000) > 20'b10000000000000000000 &&
	     dlyHoldoffBytes >= bytesWritten &&
	     dlyHoldoffCycles >= cyclesPassed ;
  assign NOT_mesgRF_rRdPtr_52_PLUS_512_93_EQ_mesgRF_rWr_ETC___d208 =
	     mesgRF_rRdPtr + 11'b01000000000 != mesgRF_rWrPtr &&
	     (!rdSerEmpty && rdSerPos != 2'b00 || wide16Fb__EMPTY_N) ;
  assign NOT_wsiS_reqFifo_countReg_96_ULE_1_97___d698 =
	     wsiS_reqFifo_countReg > 2'b01 ;
  assign _dor1bytesWritten__EN_write =
	     WILL_FIRE_RL_wmwt_messagePushPrecise ||
	     WILL_FIRE_RL_wmwt_messagePushImprecise ;
  assign addr__h20994 = { 12'b00, x__h21052 } ;
  assign addr__h21166 = { 12'b00, x__h21211 } ;
  assign mesg__h22346 = mesgRF_wDataOut__wget ;
  assign metaRF_RDY_enq__41_AND_NOT_rdSerEmpty_96_97_AN_ETC___d242 =
	     metaRF__FULL_N &&
	     (!rdSerEmpty && rdSerPos != 2'b00 || wide16Fb__EMPTY_N) ;
  assign metaWF_RDY_deq__58_AND_NOT_wrtSerPos_11_EQ_3_1_ETC___d365 =
	     metaWF__EMPTY_N &&
	     (wrtSerPos != 2'b11 && metaWF__D_OUT[23:0] != 24'b000000000000000000000000 ||
	      IF_wrtSerPos_11_EQ_0_12_OR_wrtSerPos_11_EQ_1_1_ETC___d904) ;
  assign mlp1__h17953 = MUX_mesgLengthSoFar__write_1__VAL_2 ;
  assign rdat__h21847 = { 8'b00000000, x__h21850 } ;
  assign rdat__h22030 = { 12'b00, dlyWordsStored_value } ;
  assign rdat__h22038 = { 24'b000000000000000000000000, dlyReadCredit_value } ;
  assign rdat__h22046 = { 12'b00, dlyWAG } ;
  assign rdat__h22054 = { 12'b00, dlyRAG } ;
  assign v__h22720 = metaRF__D_IN ;
  assign wci_cState_9_EQ_2_0_AND_dlyCtrl_4_BITS_3_TO_0__ETC___d397 =
	     wci_cState == 3'b010 && dlyCtrl[3:0] == 4'h7 && mesgLength[14] &&
	     !doAbort &&
	     (preciseBurst && wsiWordsRemain == 12'b00 ||
	      impreciseBurst && endOfMessage) ;
  assign wrtSerPos_11_PLUS_1___d1014 = wrtSerPos + 2'b01 ;
  assign x1__h19969 = { 96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, x__h19905[31:0] } ;
  assign x1__h19978 = { 64'b0000000000000000000000000000000000000000000000000000000000000000, x__h19905[31:0], wrtSerStage } ;
  assign x1__h20492 = { 96'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000, metaWF__D_OUT } ;
  assign x1__h20501 = { 64'b0000000000000000000000000000000000000000000000000000000000000000, metaWF__D_OUT, wrtSerStage } ;
  assign x1_length__h17254 = { 10'b0000000000, x__h17298 } ;
  assign x1_opcode__h17253 = opcode[8] ? opcode[7:0] : 8'b00000000 ;
  assign x__h15126 = mesgWF_rRdPtr + 11'b1 ;
  assign x__h15234 =
	     mesgWF_pwEnqueue__whas ? wsiS_reqFifo__D_OUT[295:40] : 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
  assign x__h16052 = mesgRF_rRdPtr + 11'b1 ;
  assign x__h16160 = CAN_FIRE_RL_rdSer_body ? mesgRF_wDataIn__wget : 256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000 ;
  assign x__h17298 = mesgLength[14] ? mesgLength[13:0] : 14'b00000000000000 ;
  assign x__h19905 = mesgWF_wDataOut__wget ;
  assign x__h21052 = { dlyRAG, 4'h0 } ;
  assign x__h21211 = { dlyWAG, 4'h0 } ;
  assign x__h21850 = { wmemi_statusR, wsiS_statusR, wsiM_statusR } ;
  assign x_burstLength__h22437 =
	     (readMeta[23:0] == 24'b000000000000000000000000) ? 12'b01 : readMeta[16:5] ;
  assign x_byteEn__h22438 = (readMeta[23:0] == 24'b000000000000000000000000) ? 32'b00000000000000000000000000000000 : 32'hFFFFFFFF ;
  always@(wci_reqF__D_OUT or
	  dlyCtrl or
	  dlyHoldoffBytes or
	  dlyHoldoffCycles or
	  mesgWtCount or
	  mesgRdCount or
	  bytesWritten or
	  rdat__h21847 or
	  wsiS_extStatusW__wget or
	  wsiM_extStatusW__wget or
	  wmemiWrReq or
	  wmemiRdReq or
	  wmemiRdResp or
	  rdat__h22030 or rdat__h22038 or rdat__h22046 or rdat__h22054)
  begin
    case (wci_reqF__D_OUT[51:32])
      20'h0: x_data__h21804 = dlyCtrl;
      20'h00004: x_data__h21804 = dlyHoldoffBytes;
      20'h00008: x_data__h21804 = dlyHoldoffCycles;
      20'h0000C: x_data__h21804 = mesgWtCount;
      20'h00010: x_data__h21804 = mesgRdCount;
      20'h00014: x_data__h21804 = bytesWritten;
      20'h00018: x_data__h21804 = rdat__h21847;
      20'h0001C: x_data__h21804 = 32'b00000000000000000000000000000000;
      20'h00020: x_data__h21804 = wsiS_extStatusW__wget[95:64];
      20'h00024: x_data__h21804 = wsiS_extStatusW__wget[63:32];
      20'h00028: x_data__h21804 = wsiS_extStatusW__wget[31:0];
      20'h0002C: x_data__h21804 = wsiM_extStatusW__wget[95:64];
      20'h00030: x_data__h21804 = wsiM_extStatusW__wget[63:32];
      20'h00034: x_data__h21804 = wsiM_extStatusW__wget[31:0];
      20'h00038: x_data__h21804 = wmemiWrReq;
      20'h0003C: x_data__h21804 = wmemiRdReq;
      20'h00040: x_data__h21804 = wmemiRdResp;
      20'h00044: x_data__h21804 = rdat__h22030;
      20'h00048: x_data__h21804 = rdat__h22038;
      20'h0004C: x_data__h21804 = rdat__h22046;
      20'h00050: x_data__h21804 = rdat__h22054;
      default: x_data__h21804 = 32'b00000000000000000000000000000000;
    endcase
  end
  always@(wrtSerPos or wide16Fa__FULL_N)
  begin
    case (wrtSerPos)
     // 2'b00, 2'b01, 2'b10
	 2'b10:
	  IF_wrtSerPos_11_EQ_0_12_OR_wrtSerPos_11_EQ_1_1_ETC___d904 =
	      wide16Fa__FULL_N;
		   2'b00:
	  IF_wrtSerPos_11_EQ_0_12_OR_wrtSerPos_11_EQ_1_1_ETC___d904 =
	      wide16Fa__FULL_N;
		   2'b01:
	  IF_wrtSerPos_11_EQ_0_12_OR_wrtSerPos_11_EQ_1_1_ETC___d904 =
	      wide16Fa__FULL_N;
      2'b11:
	  IF_wrtSerPos_11_EQ_0_12_OR_wrtSerPos_11_EQ_1_1_ETC___d904 =
	      wrtSerPos != 2'b11 || wide16Fa__FULL_N;
    endcase
  end
  always@(wrtSerPos)
  begin
    case (wrtSerPos)
     // 2'b00, 2'b01, 2'b10, 2'b11: CASE_wrtSerPos_0b1_0_1_1_1_2_1_3_0b1__q1 = 1'b1;
	 2'b00: CASE_wrtSerPos_0b1_0_1_1_1_2_1_3_0b1__q1 = 1'b1;
	 2'b01: CASE_wrtSerPos_0b1_0_1_1_1_2_1_3_0b1__q1 = 1'b1;
	 2'b10: CASE_wrtSerPos_0b1_0_1_1_1_2_1_3_0b1__q1 = 1'b1;
	 2'b11: CASE_wrtSerPos_0b1_0_1_1_1_2_1_3_0b1__q1 = 1'b1;
    endcase
  end

  // handling of inlined registers

  always@(posedge wciS0_Clk)
  begin
    if (!wciS0_MReset_n)
      begin
        abortCount <=  32'b00000000000000000000000000000000;
	blockDelayWrite <=  1'b0;
	bytesRead <=  32'b00;
	bytesWritten <=  32'b00000000000000000000000000000000;
	cyclesPassed <=  32'b00000000000000000000000000000000;
	dlyCtrl <=  dlyCtrlInit;
	dlyHoldoffBytes <=  32'b00000000000000000000000000000000;
	dlyHoldoffCycles <=  32'b00000000000000000000000000000000;
	dlyRAG <=  20'b00000000000000000000;
	dlyReadCredit_value <=  8'b00000000;
	dlyWAG <=  20'b00000000000000000000;
	dlyWordsStored_value <=  20'b00000000000000000000;
	doAbort <=  1'b0;
	endOfMessage <=  1'b0;
//	errCount <=  256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
	impreciseBurst <=  1'b0;
	mesgLength <=  15'b010101010101010;
	mesgLengthSoFar <=  14'b00000000000000;
	mesgRF_rCache <= 
	    268'h2AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
	mesgRF_rRdPtr <=  11'b0;
	mesgRF_rWrPtr <=  11'b0;
	mesgRdCount <=  32'b00000000000000000000000000000000;
	mesgReqValid <=  1'b0;
	mesgWF_rCache <= 
	    268'h2AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
	mesgWF_rRdPtr <=  11'b0;
	mesgWF_rWrPtr <=  11'b0;
	mesgWtCount <=  32'b00000000000000000000000000000000;
	opcode <=  9'b010101010;
	preciseBurst <=  1'b0;
	rdSerAddr <=  32'b00000000000000000000000000000000;
	rdSerEmpty <=  1'b1;
	rdSerPos <=  2'b00;
	rdSerUnroll <=  16'b0000000000000000;
	rdSyncWord <=  1'b0;
	readyToPush <=  1'b0;
	readyToRequest <=  1'b0;
	unrollCnt <=  16'b0000000000000000;
//	valExpect <=  256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
	wci_cEdge <=  3'b111;
	wci_cState <=  3'b000;
	wci_ctlAckReg <=  1'b0;
	wci_ctlOpActive <=  1'b0;
	wci_illegalEdge <=  1'b0;
	wci_nState <=  3'b000;
	wci_reqF_countReg <=  2'b00;
	wci_respF_c_r <=  2'b00;
	wci_respF_q_0 <=  34'h0AAAAAAAA;
	wci_respF_q_1 <=  34'h0AAAAAAAA;
	wci_sFlagReg <=  1'b0;
	wci_sThreadBusy_d <=  1'b1;
	wmemiRdReq <=  32'b00000000000000000000000000000000;
	wmemiRdResp <=  32'b00000000000000000000000000000000;
	wmemiWrReq <=  32'b00000000000000000000000000000000;
	wmemi_busyWithMessage <=  1'b0;
	wmemi_dhF_c_r <=  2'b00;
	wmemi_dhF_q_0 <= 
	    146'h0AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
	wmemi_dhF_q_1 <= 
	    146'h0AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
	wmemi_errorSticky <=  1'b0;
	wmemi_operateD <=  1'b0;
	wmemi_peerIsReady <=  1'b1;
	wmemi_reqF_c_r <=  2'b00;
	wmemi_reqF_q_0 <=  52'h0AAAAAAAAAAAA;
	wmemi_reqF_q_1 <=  52'h0AAAAAAAAAAAA;
	wmemi_trafficSticky <=  1'b0;
	wrtDutyCount <=  3'b000;
	wrtSerAddr <=  32'b00000000000000000000000000000000;
	wrtSerPos <=  2'b00;
	wrtSerUnroll <=  16'b0000000000000000;
	wsiM_burstKind <=  2'b00;
	wsiM_errorSticky <=  1'b0;
	wsiM_iMesgCount <=  32'b00000000000000000000000000000000;
	wsiM_operateD <=  1'b0;
	wsiM_pMesgCount <=  32'b00000000000000000000000000000000;
	wsiM_peerIsReady <=  1'b0;
	wsiM_reqFifo_c_r <=  2'b00;
	wsiM_reqFifo_q_0 <= 
	    313'h00000AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA00;
	wsiM_reqFifo_q_1 <= 
	    313'h00000AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA00;
	wsiM_sThreadBusy_d <=  1'b1;
	wsiM_tBusyCount <=  32'b00000000000000000000000000000000;
	wsiM_trafficSticky <=  1'b0;
	wsiS_burstKind <=  2'b00;
	wsiS_errorSticky <=  1'b0;
	wsiS_iMesgCount <=  32'b00000000000000000000000000000000;
	wsiS_operateD <=  1'b0;
	wsiS_pMesgCount <=  32'b00000000000000000000000000000000;
	wsiS_peerIsReady <=  1'b0;
	wsiS_reqFifo_countReg <=  2'b00;
	wsiS_tBusyCount <=  32'b00000000000000000000000000000000;
	wsiS_trafficSticky <=  1'b0;
	wsiWordsRemain <=  12'b00;
	zeroLengthMesg <=  1'b0;
      end
    else
      begin
        if (abortCount__EN)
	  abortCount <=  abortCount__D_IN;
	if (blockDelayWrite__EN)
	  blockDelayWrite <=  blockDelayWrite__D_IN;
	if (bytesRead__EN) bytesRead <=  bytesRead__D_IN;
	if (bytesWritten__EN)
	  bytesWritten <=  bytesWritten__D_IN;
	if (cyclesPassed__EN)
	  cyclesPassed <=  cyclesPassed__D_IN;
	if (dlyCtrl__EN) dlyCtrl <=  dlyCtrl__D_IN;
	if (dlyHoldoffBytes__EN)
	  dlyHoldoffBytes <=  dlyHoldoffBytes__D_IN;
	if (dlyHoldoffCycles__EN)
	  dlyHoldoffCycles <=  dlyHoldoffCycles__D_IN;
	if (dlyRAG__EN) dlyRAG <=  dlyRAG__D_IN;
	if (dlyReadCredit_value__EN)
	  dlyReadCredit_value <= 
	      dlyReadCredit_value__D_IN;
	if (dlyWAG__EN) dlyWAG <=  dlyWAG__D_IN;
	if (dlyWordsStored_value__EN)
	  dlyWordsStored_value <= 
	      dlyWordsStored_value__D_IN;
	if (doAbort__EN) doAbort <=  doAbort__D_IN;
	if (endOfMessage__EN)
	  endOfMessage <=  endOfMessage__D_IN;
//	if (errCount__EN) errCount <=  errCount__D_IN;
	if (impreciseBurst__EN)
	  impreciseBurst <=  impreciseBurst__D_IN;
	if (mesgLength__EN)
	  mesgLength <=  mesgLength__D_IN;
	if (mesgLengthSoFar__EN)
	  mesgLengthSoFar <=  mesgLengthSoFar__D_IN;
	if (mesgRF_rCache__EN)
	  mesgRF_rCache <=  mesgRF_rCache__D_IN;
	if (mesgRF_rRdPtr__EN)
	  mesgRF_rRdPtr <=  mesgRF_rRdPtr__D_IN;
	if (mesgRF_rWrPtr__EN)
	  mesgRF_rWrPtr <=  mesgRF_rWrPtr__D_IN;
	if (mesgRdCount__EN)
	  mesgRdCount <=  mesgRdCount__D_IN;
	if (mesgReqValid__EN)
	  mesgReqValid <=  mesgReqValid__D_IN;
	if (mesgWF_rCache__EN)
	  mesgWF_rCache <=  mesgWF_rCache__D_IN;
	if (mesgWF_rRdPtr__EN)
	  mesgWF_rRdPtr <=  mesgWF_rRdPtr__D_IN;
	if (mesgWF_rWrPtr__EN)
	  mesgWF_rWrPtr <=  mesgWF_rWrPtr__D_IN;
	if (mesgWtCount__EN)
	  mesgWtCount <=  mesgWtCount__D_IN;
	if (opcode__EN) opcode <=  opcode__D_IN;
	if (preciseBurst__EN)
	  preciseBurst <=  preciseBurst__D_IN;
	if (rdSerAddr__EN) rdSerAddr <=  rdSerAddr__D_IN;
	if (rdSerEmpty__EN)
	  rdSerEmpty <=  rdSerEmpty__D_IN;
	if (rdSerPos__EN) rdSerPos <=  rdSerPos__D_IN;
	if (rdSerUnroll__EN)
	  rdSerUnroll <=  rdSerUnroll__D_IN;
	if (rdSyncWord__EN)
	  rdSyncWord <=  rdSyncWord__D_IN;
	if (readyToPush__EN)
	  readyToPush <=  readyToPush__D_IN;
	if (readyToRequest__EN)
	  readyToRequest <=  readyToRequest__D_IN;
	if (unrollCnt__EN) unrollCnt <=  unrollCnt__D_IN;
//	if (valExpect__EN) valExpect <=  valExpect__D_IN;
	if (wci_cEdge__EN) wci_cEdge <=  wci_cEdge__D_IN;
	if (wci_cState__EN)
	  wci_cState <=  wci_cState__D_IN;
	if (wci_ctlAckReg__EN)
	  wci_ctlAckReg <=  wci_ctlAckReg__D_IN;
	if (wci_ctlOpActive__EN)
	  wci_ctlOpActive <=  wci_ctlOpActive__D_IN;
	if (wci_illegalEdge__EN)
	  wci_illegalEdge <=  wci_illegalEdge__D_IN;
	if (wci_nState__EN)
	  wci_nState <=  wci_nState__D_IN;
	if (wci_reqF_countReg__EN)
	  wci_reqF_countReg <=  wci_reqF_countReg__D_IN;
	if (wci_respF_c_r__EN)
	  wci_respF_c_r <=  wci_respF_c_r__D_IN;
	if (wci_respF_q_0__EN)
	  wci_respF_q_0 <=  wci_respF_q_0__D_IN;
	if (wci_respF_q_1__EN)
	  wci_respF_q_1 <=  wci_respF_q_1__D_IN;
	if (wci_sFlagReg__EN)
	  wci_sFlagReg <=  wci_sFlagReg__D_IN;
	if (wci_sThreadBusy_d__EN)
	  wci_sThreadBusy_d <=  wci_sThreadBusy_d__D_IN;
	if (wmemiRdReq__EN)
	  wmemiRdReq <=  wmemiRdReq__D_IN;
	if (wmemiRdResp__EN)
	  wmemiRdResp <=  wmemiRdResp__D_IN;
	if (wmemiWrReq__EN)
	  wmemiWrReq <=  wmemiWrReq__D_IN;
	if (wmemi_busyWithMessage__EN)
	  wmemi_busyWithMessage <= 
	      wmemi_busyWithMessage__D_IN;
	if (wmemi_dhF_c_r__EN)
	  wmemi_dhF_c_r <=  wmemi_dhF_c_r__D_IN;
	if (wmemi_dhF_q_0__EN)
	  wmemi_dhF_q_0 <=  wmemi_dhF_q_0__D_IN;
	if (wmemi_dhF_q_1__EN)
	  wmemi_dhF_q_1 <=  wmemi_dhF_q_1__D_IN;
	if (wmemi_errorSticky__EN)
	  wmemi_errorSticky <=  wmemi_errorSticky__D_IN;
	if (wmemi_operateD__EN)
	  wmemi_operateD <=  wmemi_operateD__D_IN;
	if (wmemi_peerIsReady__EN)
	  wmemi_peerIsReady <=  wmemi_peerIsReady__D_IN;
	if (wmemi_reqF_c_r__EN)
	  wmemi_reqF_c_r <=  wmemi_reqF_c_r__D_IN;
	if (wmemi_reqF_q_0__EN)
	  wmemi_reqF_q_0 <=  wmemi_reqF_q_0__D_IN;
	if (wmemi_reqF_q_1__EN)
	  wmemi_reqF_q_1 <=  wmemi_reqF_q_1__D_IN;
	if (wmemi_trafficSticky__EN)
	  wmemi_trafficSticky <= 
	      wmemi_trafficSticky__D_IN;
	if (wrtDutyCount__EN)
	  wrtDutyCount <=  wrtDutyCount__D_IN;
	if (wrtSerAddr__EN)
	  wrtSerAddr <=  wrtSerAddr__D_IN;
	if (wrtSerPos__EN) wrtSerPos <=  wrtSerPos__D_IN;
	if (wrtSerUnroll__EN)
	  wrtSerUnroll <=  wrtSerUnroll__D_IN;
	if (wsiM_burstKind__EN)
	  wsiM_burstKind <=  wsiM_burstKind__D_IN;
	if (wsiM_errorSticky__EN)
	  wsiM_errorSticky <=  wsiM_errorSticky__D_IN;
	if (wsiM_iMesgCount__EN)
	  wsiM_iMesgCount <=  wsiM_iMesgCount__D_IN;
	if (wsiM_operateD__EN)
	  wsiM_operateD <=  wsiM_operateD__D_IN;
	if (wsiM_pMesgCount__EN)
	  wsiM_pMesgCount <=  wsiM_pMesgCount__D_IN;
	if (wsiM_peerIsReady__EN)
	  wsiM_peerIsReady <=  wsiM_peerIsReady__D_IN;
	if (wsiM_reqFifo_c_r__EN)
	  wsiM_reqFifo_c_r <=  wsiM_reqFifo_c_r__D_IN;
	if (wsiM_reqFifo_q_0__EN)
	  wsiM_reqFifo_q_0 <=  wsiM_reqFifo_q_0__D_IN;
	if (wsiM_reqFifo_q_1__EN)
	  wsiM_reqFifo_q_1 <=  wsiM_reqFifo_q_1__D_IN;
	if (wsiM_sThreadBusy_d__EN)
	  wsiM_sThreadBusy_d <=  wsiM_sThreadBusy_d__D_IN;
	if (wsiM_tBusyCount__EN)
	  wsiM_tBusyCount <=  wsiM_tBusyCount__D_IN;
	if (wsiM_trafficSticky__EN)
	  wsiM_trafficSticky <=  wsiM_trafficSticky__D_IN;
	if (wsiS_burstKind__EN)
	  wsiS_burstKind <=  wsiS_burstKind__D_IN;
	if (wsiS_errorSticky__EN)
	  wsiS_errorSticky <=  wsiS_errorSticky__D_IN;
	if (wsiS_iMesgCount__EN)
	  wsiS_iMesgCount <=  wsiS_iMesgCount__D_IN;
	if (wsiS_operateD__EN)
	  wsiS_operateD <=  wsiS_operateD__D_IN;
	if (wsiS_pMesgCount__EN)
	  wsiS_pMesgCount <=  wsiS_pMesgCount__D_IN;
	if (wsiS_peerIsReady__EN)
	  wsiS_peerIsReady <=  wsiS_peerIsReady__D_IN;
	if (wsiS_reqFifo_countReg__EN)
	  wsiS_reqFifo_countReg <= 
	      wsiS_reqFifo_countReg__D_IN;
	if (wsiS_tBusyCount__EN)
	  wsiS_tBusyCount <=  wsiS_tBusyCount__D_IN;
	if (wsiS_trafficSticky__EN)
	  wsiS_trafficSticky <=  wsiS_trafficSticky__D_IN;
	if (wsiWordsRemain__EN)
	  wsiWordsRemain <=  wsiWordsRemain__D_IN;
	if (zeroLengthMesg__EN)
	  zeroLengthMesg <=  zeroLengthMesg__D_IN;
      end
    if (rdSerMeta__EN) rdSerMeta <=  rdSerMeta__D_IN;
    if (rdSerStage__EN) rdSerStage <=  rdSerStage__D_IN;
    if (rdSerStage_1__EN)
      rdSerStage_1 <=  rdSerStage_1__D_IN;
    if (rdSerStage_2__EN)
      rdSerStage_2 <=  rdSerStage_2__D_IN;
    if (rdSerStage_3__EN)
      rdSerStage_3 <=  rdSerStage_3__D_IN;
    if (readMeta__EN) readMeta <=  readMeta__D_IN;
    if (wmemi_statusR__EN)
      wmemi_statusR <=  wmemi_statusR__D_IN;
    if (wrtSerMeta__EN) wrtSerMeta <=  wrtSerMeta__D_IN;
    if (wrtSerStage__EN) wrtSerStage <=  wrtSerStage__D_IN;
    if (wrtSerStage_1__EN)
      wrtSerStage_1 <=  wrtSerStage_1__D_IN;
    if (wrtSerStage_2__EN)
      wrtSerStage_2 <=  wrtSerStage_2__D_IN;
    if (wrtSerStage_3__EN)
      wrtSerStage_3 <=  wrtSerStage_3__D_IN;
    if (wsiM_statusR__EN)
      wsiM_statusR <=  wsiM_statusR__D_IN;
    if (wsiS_statusR__EN)
      wsiS_statusR <=  wsiS_statusR__D_IN;
  end

  // handling of system tasks


endmodule  // mkDelayWorker32B


 
 
module ResetToBool (RST, VAL);

input RST;
output VAL;
reg VAL;

always @ (RST or VAL)
begin

if (RST == 1)
VAL=1'b0;

end
endmodule

 
module arSRLFIFO_a (CLK, RST_N, D_IN,ENQ,DEQ,CLR,D_OUT,EMPTY_N,FULL_N);

input CLK;
input RST_N;
input [31:0] D_IN;
input ENQ;
input DEQ;
input CLR;
output [31:0] D_OUT;
output EMPTY_N;
output FULL_N;



wire fulln;
wire emptyn;

wire always_one;
wire always_zero;

assign always_one = 1'b1;
assign always_zero = 1'b0;

generic_fifo_sc_a fifo_1
(.clk(CLK),
 .rst(RST_N),
 .clr (CLR),
 .din (D_IN),
 .we (ENQ),
 .dout (D_OUT),
 .re (DEQ),
 .full_r (FULL_N),
 .empty_r(EMPTY_N),
 .full_n_r (fulln),
 .empty_n_r (emptyn)
 );
 







endmodule








/////////////////////////////////////////////////////////////////////
////                                                             ////
////  Universal FIFO Single Clock                                ////
////                                                             ////
////                                                             ////
////  Author: Rudolf Usselmann                                   ////
////          rudi@asics.ws                                      ////
////                                                             ////
////                                                             ////
////  D/L from: http://www.opencores.org/cores/generic_fifos/    ////
////                                                             ////
/////////////////////////////////////////////////////////////////////
////                                                             ////
//// Copyright (C) 2000-2002 Rudolf Usselmann                    ////
////                         www.asics.ws                        ////
////                         rudi@asics.ws                       ////
////                                                             ////
//// This source file may be used and distributed without        ////
//// restriction provided that this copyright statement is not   ////
//// removed from the file and that any derivative work contains ////
//// the original copyright notice and the associated disclaimer.////
////                                                             ////
////     THIS SOFTWARE IS PROVIDED ``AS IS'' AND WITHOUT ANY     ////
//// EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED   ////
//// TO, THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS   ////
//// FOR A PARTICULAR PURPOSE. IN NO EVENT SHALL THE AUTHOR      ////
//// OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT, INDIRECT,         ////
//// INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES    ////
//// (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE   ////
//// GOODS OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR        ////
//// BUSINESS INTERRUPTION) HOWEVER CAUSED AND ON ANY THEORY OF  ////
//// LIABILITY, WHETHER IN  CONTRACT, STRICT LIABILITY, OR TORT  ////
//// (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT  ////
//// OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED OF THE         ////
//// POSSIBILITY OF SUCH DAMAGE.                                 ////
////                                                             ////
/////////////////////////////////////////////////////////////////////
 
//  CVS Log
//
//  __Id: generic_fifo_sc_a.v,v 1.1.1.1 2002-09-25 05:42:06 rudi Exp __
//
//  __Date: 2002-09-25 05:42:06 __
//  __Revision: 1.1.1.1 __
//  __Author: rudi __
//  __Locker:  __
//  __State: Exp __
//
// Change History:
//               __Log: not supported by cvs2svn __
//
//
//
//
//
//
//
//
//
//
 
 
/*
 
Description
===========
 
I/Os
----
rst	low active, either sync. or async. master reset (see below how to select)
clr	synchronous clear (just like reset but always synchronous), high active
re	read enable, synchronous, high active
we	read enable, synchronous, high active
din	Data Input
dout	Data Output
 
full	Indicates the FIFO is full (combinatorial output)
full_r	same as above, but registered output (see note below)
empty	Indicates the FIFO is empty
empty_r	same as above, but registered output (see note below)
 
full_n		Indicates if the FIFO has space for N entries (combinatorial output)
full_n_r	same as above, but registered output (see note below)
empty_n		Indicates the FIFO has at least N entries (combinatorial output)
empty_n_r	same as above, but registered output (see note below)
 
level		indicates the FIFO level:
		2'b00	0-25%	 full
		2'b01	25-50%	 full
		2'b10	50-75%	 full
		2'b11	%75-100% full
 
combinatorial vs. registered status outputs
-------------------------------------------
Both the combinatorial and registered status outputs have exactly the same
synchronous timing. Meaning they are being asserted immediately at the clock
edge after the last read or write. The combinatorial outputs however, pass
through several levels of logic before they are output. The registered status
outputs are direct outputs of a flip-flop. The reason both are provided, is
that the registered outputs require quite a bit of additional logic inside
the FIFO. If you can meet timing of your device with the combinatorial
outputs, use them ! The FIFO will be smaller. If the status signals are
in the critical pass, use the registered outputs, they have a much smaller
output delay (actually only Tcq).
 
Parameters
----------
The FIFO takes 3 parameters:
dw	Data bus width
aw	Address bus width (Determines the FIFO size by evaluating 2^aw)
n	N is a second status threshold constant for full_n and empty_n
	If you have no need for the second status threshold, do not
	connect the outputs and the logic should be removed by your
	synthesis tool.
 
Synthesis Results
-----------------
In a Spartan 2e a 8 bit wide, 8 entries deep FIFO, takes 85 LUTs and runs
at about 116 MHz (IO insertion disabled). The registered status outputs
are valid after 2.1NS, the combinatorial once take out to 6.5 NS to be
available.
 
 
Misc
----
This design assumes you will do appropriate status checking externally.
 
IMPORTANT ! writing while the FIFO is full or reading while the FIFO is
empty will place the FIFO in an undefined state.
 
*/
 
 
// Selecting Sync. or Async Reset
// ------------------------------
// Uncomment one of the two lines below. The first line for
// synchronous reset, the second for asynchronous reset
 
//`define SC_FIFO_ASYNC_RESET				// Uncomment for Syncr. reset
//`define SC_FIFO_ASYNC_RESET	or negedge rst		// Uncomment for Async. reset

/*
parameter dw=8;
parameter aw=8;
parameter n=32;
parameter max_size = 1<<aw;
 */
 
 `define dwa 32
 `define awa 4
 
module generic_fifo_sc_a(clk, rst, clr, din, we, dout, re,
			 full_r, empty_r,
			 full_n_r, empty_n_r);
 /*
parameter dw=8;
parameter aw=8;
parameter n=32;
parameter max_size = 1<<aw;
 */
input			clk, rst, clr;
input	[`dwa-1:0]	din;
input			we;
output	[`dwa-1:0]	dout;
input			re;
wire			full; output full_r;
wire			empty; output empty_r;
wire			full_n; output full_n_r;
wire			empty_n; output empty_n_r;
wire	[1:0]		level;
 
////////////////////////////////////////////////////////////////////
//
// Local Wires
//
 
reg	[`awa-1:0]	wp;
wire	[`awa-1:0]	wp_pl1;
wire	[`awa-1:0]	wp_pl2;
reg	[`awa-1:0]	rp;
wire	[`awa-1:0]	rp_pl1;
reg			full_r;
reg			empty_r;
reg			gb;
reg			gb2;
reg	[`awa:0]		cnt;
wire			full_n, empty_n;
reg			full_n_r, empty_n_r;
 
////////////////////////////////////////////////////////////////////
//
// Memory Block
//
 wire always_zero;
 assign always_zero = 1'b0;
 wire [`dwa-1:0] junk_out;
 
 wire [`dwa-1:0] junk_in;
 
 // manually assign
 assign junk_in = 32'b00000000000000000000000000000000;
 
 // aryap: removed for benchmark
dual_port_ram #( .ADDR_WIDTH(4), .DATA_WIDTH(32))   ram1(
	.clk(		clk		),
	.addr1(		rp		),
	.addr2(		wp		),
	.we1(		we		),
	.we2(		always_zero		),
	.out1(		dout		),
	.out2(		junk_out		),
	.data1(		din		),
	.data2 (	junk_in)
	);
 
////////////////////////////////////////////////////////////////////
//
// Misc Logic
//
 
always @(posedge clk )
	if(!rst)	wp <=  {4'b0000};
	else
	if(clr)		wp <=  {4'b0000};
	else
	if(we)		wp <=  wp_pl1;
 
assign wp_pl1 = wp + { {3'b000}, 1'b1};
assign wp_pl2 = wp + { {2'b00}, 2'b10};
 
always @(posedge clk )
	if(!rst)	rp <=  {4'b0000};
	else
	if(clr)		rp <=  {4'b0000};
	else
	if(re)		rp <=  rp_pl1;
 
assign rp_pl1 = rp + { {3'b000}, 1'b1};
 
////////////////////////////////////////////////////////////////////
//
// Combinatorial Full & Empty Flags
//
 
assign empty = ((wp == rp) & !gb);
assign full  = ((wp == rp) &  gb);
 
// Guard Bit ...
always @(posedge clk )
	if(!rst)			gb <=  1'b0;
	else
	if(clr)				gb <=  1'b0;
	else
	if((wp_pl1 == rp) & we)		gb <=  1'b1;
	else
	if(re)				gb <=  1'b0;
 
////////////////////////////////////////////////////////////////////
//
// Registered Full & Empty Flags
//
 
// Guard Bit ...
always @(posedge clk )
	if(!rst)			gb2 <=  1'b0;
	else
	if(clr)				gb2 <=  1'b0;
	else
	if((wp_pl2 == rp) & we)		gb2 <=  1'b1;
	else
	if((wp != rp) & re)		gb2 <=  1'b0;
 
always @(posedge clk )
	if(!rst)				full_r <=  1'b0;
	else
	if(clr)					full_r <=  1'b0;
	else
	if(we & ((wp_pl1 == rp) & gb2) & !re)	full_r <=  1'b1;
	else
	if(re & ((wp_pl1 != rp) | !gb2) & !we)	full_r <=  1'b0;
 
always @(posedge clk )
	if(!rst)				empty_r <=  1'b1;
	else
	if(clr)					empty_r <=  1'b1;
	else
	if(we & ((wp != rp_pl1) | gb2) & !re)	empty_r <=  1'b0;
	else
	if(re & ((wp == rp_pl1) & !gb2) & !we)	empty_r <=  1'b1;
 
////////////////////////////////////////////////////////////////////
//
// Combinatorial Full_n & Empty_n Flags
//
 
assign empty_n = cnt < `n;
assign full_n  = !(cnt < (`max_size-`n+1));
assign level = {{cnt[`awa]}, {cnt[`awa]}} | cnt[`awa-1:`awa-2];
 
// N entries status
always @(posedge clk )
	if(!rst)	cnt <=  {4'b0000};
	else
	if(clr)		cnt <=  {4'b0000};
	else
	if( re & !we)	cnt <=  cnt + { 5'b11111};
	else
	if(!re &  we)	cnt <=  cnt + { {4'b0000}, 1'b1};
 
////////////////////////////////////////////////////////////////////
//
// Registered Full_n & Empty_n Flags
//
 
always @(posedge clk )
	if(!rst)				empty_n_r <=  1'b1;
	else
	if(clr)					empty_n_r <=  1'b1;
	else
	if(we & (cnt >= (`n-1) ) & !re)		empty_n_r <=  1'b0;
	else
	if(re & (cnt <= `n ) & !we)		empty_n_r <=  1'b1;
 
always @(posedge clk )
	if(!rst)				full_n_r <=  1'b0;
	else
	if(clr)					full_n_r <=  1'b0;
	else
	if(we & (cnt >= (`max_size-`n) ) & !re)	full_n_r <=  1'b1;
	else
	if(re & (cnt <= (`max_size-`n+1)) & !we)	full_n_r <=  1'b0;

endmodule
 

module arSRLFIFO_b (CLK, RST_N, D_IN,ENQ,DEQ,CLR,D_OUT,EMPTY_N,FULL_N);

input CLK;
input RST_N;
input [31:0] D_IN;
input ENQ;
input DEQ;
input CLR;
output [31:0] D_OUT;
output EMPTY_N;
output FULL_N;



wire fulln;
wire emptyn;

wire always_one;
wire always_zero;

assign always_one = 1'b1;
assign always_zero = 1'b0;

generic_fifo_sc_b fifo_1
(.clk(CLK),
 .rst(RST_N),
 .clr (CLR),
 .din (D_IN),
 .we (ENQ),
 .dout (D_OUT),
 .re (DEQ),
 .full_r (FULL_N),
 .empty_r(EMPTY_N),
 .full_n_r (fulln),
 .empty_n_r (emptyn)
 );
 







endmodule








/////////////////////////////////////////////////////////////////////
////                                                             ////
////  Universal FIFO Single Clock                                ////
////                                                             ////
////                                                             ////
////  Author: Rudolf Usselmann                                   ////
////          rudi@asics.ws                                      ////
////                                                             ////
////                                                             ////
////  D/L from: http://www.opencores.org/cores/generic_fifos/    ////
////                                                             ////
/////////////////////////////////////////////////////////////////////
////                                                             ////
//// Copyright (C) 2000-2002 Rudolf Usselmann                    ////
////                         www.asics.ws                        ////
////                         rudi@asics.ws                       ////
////                                                             ////
//// This source file may be used and distributed without        ////
//// restriction provided that this copyright statement is not   ////
//// removed from the file and that any derivative work contains ////
//// the original copyright notice and the associated disclaimer.////
////                                                             ////
////     THIS SOFTWARE IS PROVIDED ``AS IS'' AND WITHOUT ANY     ////
//// EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED   ////
//// TO, THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS   ////
//// FOR A PARTICULAR PURPOSE. IN NO EVENT SHALL THE AUTHOR      ////
//// OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT, INDIRECT,         ////
//// INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES    ////
//// (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE   ////
//// GOODS OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR        ////
//// BUSINESS INTERRUPTION) HOWEVER CAUSED AND ON ANY THEORY OF  ////
//// LIABILITY, WHETHER IN  CONTRACT, STRICT LIABILITY, OR TORT  ////
//// (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT  ////
//// OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED OF THE         ////
//// POSSIBILITY OF SUCH DAMAGE.                                 ////
////                                                             ////
/////////////////////////////////////////////////////////////////////
 
//  CVS Log
//
//  __Id: generic_fifo_sc_a.v,v 1.1.1.1 2002-09-25 05:42:06 rudi Exp __
//
//  __Date: 2002-09-25 05:42:06 __
//  __Revision: 1.1.1.1 __
//  __Author: rudi __
//  __Locker:  __
//  __State: Exp __
//
// Change History:
//               __Log: not supported by cvs2svn __
//
//
//
//
//
//
//
//
//
//
 
 
/*
 
Description
===========
 
I/Os
----
rst	low active, either sync. or async. master reset (see below how to select)
clr	synchronous clear (just like reset but always synchronous), high active
re	read enable, synchronous, high active
we	read enable, synchronous, high active
din	Data Input
dout	Data Output
 
full	Indicates the FIFO is full (combinatorial output)
full_r	same as above, but registered output (see note below)
empty	Indicates the FIFO is empty
empty_r	same as above, but registered output (see note below)
 
full_n		Indicates if the FIFO has space for N entries (combinatorial output)
full_n_r	same as above, but registered output (see note below)
empty_n		Indicates the FIFO has at least N entries (combinatorial output)
empty_n_r	same as above, but registered output (see note below)
 
level		indicates the FIFO level:
		2'b00	0-25%	 full
		2'b01	25-50%	 full
		2'b10	50-75%	 full
		2'b11	%75-100% full
 
combinatorial vs. registered status outputs
-------------------------------------------
Both the combinatorial and registered status outputs have exactly the same
synchronous timing. Meaning they are being asserted immediately at the clock
edge after the last read or write. The combinatorial outputs however, pass
through several levels of logic before they are output. The registered status
outputs are direct outputs of a flip-flop. The reason both are provided, is
that the registered outputs require quite a bit of additional logic inside
the FIFO. If you can meet timing of your device with the combinatorial
outputs, use them ! The FIFO will be smaller. If the status signals are
in the critical pass, use the registered outputs, they have a much smaller
output delay (actually only Tcq).
 
Parameters
----------
The FIFO takes 3 parameters:
dw	Data bus width
aw	Address bus width (Determines the FIFO size by evaluating 2^aw)
n	N is a second status threshold constant for full_n and empty_n
	If you have no need for the second status threshold, do not
	connect the outputs and the logic should be removed by your
	synthesis tool.
 
Synthesis Results
-----------------
In a Spartan 2e a 8 bit wide, 8 entries deep FIFO, takes 85 LUTs and runs
at about 116 MHz (IO insertion disabled). The registered status outputs
are valid after 2.1NS, the combinatorial once take out to 6.5 NS to be
available.
 
 
Misc
----
This design assumes you will do appropriate status checking externally.
 
IMPORTANT ! writing while the FIFO is full or reading while the FIFO is
empty will place the FIFO in an undefined state.
 
*/
 
 
// Selecting Sync. or Async Reset
// ------------------------------
// Uncomment one of the two lines below. The first line for
// synchronous reset, the second for asynchronous reset
 
//`define SC_FIFO_ASYNC_RESET				// Uncomment for Syncr. reset
//`define SC_FIFO_ASYNC_RESET	or negedge rst		// Uncomment for Async. reset

/*
parameter dw=8;
parameter aw=8;
parameter n=32;
parameter max_size = 1<<aw;
 */

 
module generic_fifo_sc_b(clk, rst, clr, din, we, dout, re,
			 full_r, empty_r,
			 full_n_r, empty_n_r);
 /*
parameter dw=8;
parameter aw=8;
parameter n=32;
parameter max_size = 1<<aw;
 */
input			clk, rst, clr;
input	[`dwa-1:0]	din;
input			we;
output	[`dwa-1:0]	dout;
input			re;
wire			full; output full_r;
wire			empty; output empty_r;
wire			full_n; output full_n_r;
wire			empty_n; output empty_n_r;
wire	[1:0]		level;
 
////////////////////////////////////////////////////////////////////
//
// Local Wires
//
 
reg	[`awa-1:0]	wp;
wire	[`awa-1:0]	wp_pl1;
wire	[`awa-1:0]	wp_pl2;
reg	[`awa-1:0]	rp;
wire	[`awa-1:0]	rp_pl1;
reg			full_r;
reg			empty_r;
reg			gb;
reg			gb2;
reg	[`awa:0]		cnt;
wire			full_n, empty_n;
reg			full_n_r, empty_n_r;
 
////////////////////////////////////////////////////////////////////
//
// Memory Block
//
 wire always_zero;
 assign always_zero = 1'b0;
 wire [`dwa-1:0] junk_out;
 
 wire [`dwa-1:0] junk_in;
 
 // manually assign
 assign junk_in = 32'b00000000000000000000000000000000;
 
 // aryap: removed for benchmark
dual_port_ram #( .ADDR_WIDTH(4), .DATA_WIDTH(32))   ram1(
	.clk(		clk		),
	.addr1(		rp		),
	.addr2(		wp		),
	.we1(		we		),
	.we2(		always_zero		),
	.out1(		dout		),
	.out2(		junk_out		),
	.data1(		din		),
	.data2 (	junk_in)
	);
 
////////////////////////////////////////////////////////////////////
//
// Misc Logic
//
 
always @(posedge clk )
	if(!rst)	wp <=  {4'b0000};
	else
	if(clr)		wp <=  {4'b0000};
	else
	if(we)		wp <=  wp_pl1;
 
assign wp_pl1 = wp + { {3'b000}, 1'b1};
assign wp_pl2 = wp + { {2'b00}, 2'b10};
 
always @(posedge clk )
	if(!rst)	rp <=  {4'b0000};
	else
	if(clr)		rp <=  {4'b0000};
	else
	if(re)		rp <=  rp_pl1;
 
assign rp_pl1 = rp + { {3'b000}, 1'b1};
 
////////////////////////////////////////////////////////////////////
//
// Combinatorial Full & Empty Flags
//
 
assign empty = ((wp == rp) & !gb);
assign full  = ((wp == rp) &  gb);
 
// Guard Bit ...
always @(posedge clk )
	if(!rst)			gb <=  1'b0;
	else
	if(clr)				gb <=  1'b0;
	else
	if((wp_pl1 == rp) & we)		gb <=  1'b1;
	else
	if(re)				gb <=  1'b0;
 
////////////////////////////////////////////////////////////////////
//
// Registered Full & Empty Flags
//
 
// Guard Bit ...
always @(posedge clk )
	if(!rst)			gb2 <=  1'b0;
	else
	if(clr)				gb2 <=  1'b0;
	else
	if((wp_pl2 == rp) & we)		gb2 <=  1'b1;
	else
	if((wp != rp) & re)		gb2 <=  1'b0;
 
always @(posedge clk )
	if(!rst)				full_r <=  1'b0;
	else
	if(clr)					full_r <=  1'b0;
	else
	if(we & ((wp_pl1 == rp) & gb2) & !re)	full_r <=  1'b1;
	else
	if(re & ((wp_pl1 != rp) | !gb2) & !we)	full_r <=  1'b0;
 
always @(posedge clk )
	if(!rst)				empty_r <=  1'b1;
	else
	if(clr)					empty_r <=  1'b1;
	else
	if(we & ((wp != rp_pl1) | gb2) & !re)	empty_r <=  1'b0;
	else
	if(re & ((wp == rp_pl1) & !gb2) & !we)	empty_r <=  1'b1;
 
////////////////////////////////////////////////////////////////////
//
// Combinatorial Full_n & Empty_n Flags
//
 
assign empty_n = cnt < `n;
assign full_n  = !(cnt < (`max_size-`n+1));
assign level = {{cnt[`awa]}, {cnt[`awa]}} | cnt[`awa-1:`awa-2];
 
// N entries status
always @(posedge clk )
	if(!rst)	cnt <=  {4'b0000};
	else
	if(clr)		cnt <=  {4'b0000};
	else
	if( re & !we)	cnt <=  cnt + { 5'b11111};
	else
	if(!re &  we)	cnt <=  cnt + { {4'b0000}, 1'b1};
 
////////////////////////////////////////////////////////////////////
//
// Registered Full_n & Empty_n Flags
//
 
always @(posedge clk )
	if(!rst)				empty_n_r <=  1'b1;
	else
	if(clr)					empty_n_r <=  1'b1;
	else
	if(we & (cnt >= (`n-1) ) & !re)		empty_n_r <=  1'b0;
	else
	if(re & (cnt <= `n ) & !we)		empty_n_r <=  1'b1;
 
always @(posedge clk )
	if(!rst)				full_n_r <=  1'b0;
	else
	if(clr)					full_n_r <=  1'b0;
	else
	if(we & (cnt >= (`max_size-`n) ) & !re)	full_n_r <=  1'b1;
	else
	if(re & (cnt <= (`max_size-`n+1)) & !we)	full_n_r <=  1'b0;

endmodule
 

 
 
module arSRLFIFO_c (CLK, RST_N, D_IN,ENQ,DEQ,CLR,D_OUT,EMPTY_N,FULL_N);

input CLK;
input RST_N;
input [127:0] D_IN;
input ENQ;
input DEQ;
input CLR;
output [127:0] D_OUT;
output EMPTY_N;
output FULL_N;



wire fulln;
wire emptyn;

wire always_one;
wire always_zero;

assign always_one = 1'b1;
assign always_zero = 1'b0;

generic_fifo_sc_c fifo_1
(.clk(CLK),
 .rst(RST_N),
 .clr (CLR),
 .din (D_IN),
 .we (ENQ),
 .dout (D_OUT),
 .re (DEQ),
 .full_r (FULL_N),
 .empty_r(EMPTY_N),
 .full_n_r (fulln),
 .empty_n_r (emptyn)
 );
 







endmodule








/////////////////////////////////////////////////////////////////////
////                                                             ////
////  Universal FIFO Single Clock                                ////
////                                                             ////
////                                                             ////
////  Author: Rudolf Usselmann                                   ////
////          rudi@asics.ws                                      ////
////                                                             ////
////                                                             ////
////  D/L from: http://www.opencores.org/cores/generic_fifos/    ////
////                                                             ////
/////////////////////////////////////////////////////////////////////
////                                                             ////
//// Copyright (C) 2000-2002 Rudolf Usselmann                    ////
////                         www.asics.ws                        ////
////                         rudi@asics.ws                       ////
////                                                             ////
//// This source file may be used and distributed without        ////
//// restriction provided that this copyright statement is not   ////
//// removed from the file and that any derivative work contains ////
//// the original copyright notice and the associated disclaimer.////
////                                                             ////
////     THIS SOFTWARE IS PROVIDED ``AS IS'' AND WITHOUT ANY     ////
//// EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED   ////
//// TO, THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS   ////
//// FOR A PARTICULAR PURPOSE. IN NO EVENT SHALL THE AUTHOR      ////
//// OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT, INDIRECT,         ////
//// INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES    ////
//// (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE   ////
//// GOODS OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR        ////
//// BUSINESS INTERRUPTION) HOWEVER CAUSED AND ON ANY THEORY OF  ////
//// LIABILITY, WHETHER IN  CONTRACT, STRICT LIABILITY, OR TORT  ////
//// (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT  ////
//// OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED OF THE         ////
//// POSSIBILITY OF SUCH DAMAGE.                                 ////
////                                                             ////
/////////////////////////////////////////////////////////////////////
 
//  CVS Log
//
//  __Id: generic_fifo_sc_a.v,v 1.1.1.1 2002-09-25 05:42:06 rudi Exp __
//
//  __Date: 2002-09-25 05:42:06 __
//  __Revision: 1.1.1.1 __
//  __Author: rudi __
//  __Locker:  __
//  __State: Exp __
//
// Change History:
//               __Log: not supported by cvs2svn __
//
//
//
//
//
//
//
//
//
//
 
 
/*
 
Description
===========
 
I/Os
----
rst	low active, either sync. or async. master reset (see below how to select)
clr	synchronous clear (just like reset but always synchronous), high active
re	read enable, synchronous, high active
we	read enable, synchronous, high active
din	Data Input
dout	Data Output
 
full	Indicates the FIFO is full (combinatorial output)
full_r	same as above, but registered output (see note below)
empty	Indicates the FIFO is empty
empty_r	same as above, but registered output (see note below)
 
full_n		Indicates if the FIFO has space for N entries (combinatorial output)
full_n_r	same as above, but registered output (see note below)
empty_n		Indicates the FIFO has at least N entries (combinatorial output)
empty_n_r	same as above, but registered output (see note below)
 
level		indicates the FIFO level:
		2'b00	0-25%	 full
		2'b01	25-50%	 full
		2'b10	50-75%	 full
		2'b11	%75-100% full
 
combinatorial vs. registered status outputs
-------------------------------------------
Both the combinatorial and registered status outputs have exactly the same
synchronous timing. Meaning they are being asserted immediately at the clock
edge after the last read or write. The combinatorial outputs however, pass
through several levels of logic before they are output. The registered status
outputs are direct outputs of a flip-flop. The reason both are provided, is
that the registered outputs require quite a bit of additional logic inside
the FIFO. If you can meet timing of your device with the combinatorial
outputs, use them ! The FIFO will be smaller. If the status signals are
in the critical pass, use the registered outputs, they have a much smaller
output delay (actually only Tcq).
 
Parameters
----------
The FIFO takes 3 parameters:
dw	Data bus width
aw	Address bus width (Determines the FIFO size by evaluating 2^aw)
n	N is a second status threshold constant for full_n and empty_n
	If you have no need for the second status threshold, do not
	connect the outputs and the logic should be removed by your
	synthesis tool.
 
Synthesis Results
-----------------
In a Spartan 2e a 8 bit wide, 8 entries deep FIFO, takes 85 LUTs and runs
at about 116 MHz (IO insertion disabled). The registered status outputs
are valid after 2.1NS, the combinatorial once take out to 6.5 NS to be
available.
 
 
Misc
----
This design assumes you will do appropriate status checking externally.
 
IMPORTANT ! writing while the FIFO is full or reading while the FIFO is
empty will place the FIFO in an undefined state.
 
*/
 
 
// Selecting Sync. or Async Reset
// ------------------------------
// Uncomment one of the two lines below. The first line for
// synchronous reset, the second for asynchronous reset
 
//`define SC_FIFO_ASYNC_RESET				// Uncomment for Syncr. reset
//`define SC_FIFO_ASYNC_RESET	or negedge rst		// Uncomment for Async. reset

/*
parameter dw=8;
parameter aw=8;
parameter n=32;
parameter max_size = 1<<aw;
 */
 
 `define dwc 128
 `define awa 4
 
module generic_fifo_sc_c(clk, rst, clr, din, we, dout, re,
			 full_r, empty_r,
			 full_n_r, empty_n_r);
 /*
parameter dw=8;
parameter aw=8;
parameter n=32;
parameter max_size = 1<<aw;
 */
input			clk, rst, clr;
input	[`dwc-1:0]	din;
input			we;
output	[`dwc-1:0]	dout;
input			re;
wire			full; output full_r;
wire			empty; output empty_r;
wire			full_n; output full_n_r;
wire			empty_n; output empty_n_r;
wire	[1:0]		level;
 
////////////////////////////////////////////////////////////////////
//
// Local Wires
//
 
reg	[`awa-1:0]	wp;
wire	[`awa-1:0]	wp_pl1;
wire	[`awa-1:0]	wp_pl2;
reg	[`awa-1:0]	rp;
wire	[`awa-1:0]	rp_pl1;
reg			full_r;
reg			empty_r;
reg			gb;
reg			gb2;
reg	[`awa:0]		cnt;
wire			full_n, empty_n;
reg			full_n_r, empty_n_r;
 
////////////////////////////////////////////////////////////////////
//
// Memory Block
//
 wire always_zero;
 assign always_zero = 1'b0;
 wire [`dwc-1:0] junk_out;
 
 wire [`dwc-1:0] junk_in;
 
 // manually assign
 assign junk_in = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
 
dual_port_ram  #( .ADDR_WIDTH(4), .DATA_WIDTH(128))  ram1(
	.clk(		clk		),
	.addr1(		rp		),
	.addr2(		wp		),
	.we1(		we		),
	.we2(		always_zero		),
	.out1(		dout		),
	.out2(		junk_out		),
	.data1(		din		),
	.data2 (	junk_in)
	);
 
////////////////////////////////////////////////////////////////////
//
// Misc Logic
//
 
always @(posedge clk )
	if(!rst)	wp <=  {4'b0000};
	else
	if(clr)		wp <=  {4'b0000};
	else
	if(we)		wp <=  wp_pl1;
 
assign wp_pl1 = wp + { {3'b000}, 1'b1};
assign wp_pl2 = wp + { {2'b00}, 2'b10};
 
always @(posedge clk )
	if(!rst)	rp <=  {4'b0000};
	else
	if(clr)		rp <=  {4'b0000};
	else
	if(re)		rp <=  rp_pl1;
 
assign rp_pl1 = rp + { {3'b000}, 1'b1};
 
////////////////////////////////////////////////////////////////////
//
// Combinatorial Full & Empty Flags
//
 
assign empty = ((wp == rp) & !gb);
assign full  = ((wp == rp) &  gb);
 
// Guard Bit ...
always @(posedge clk )
	if(!rst)			gb <=  1'b0;
	else
	if(clr)				gb <=  1'b0;
	else
	if((wp_pl1 == rp) & we)		gb <=  1'b1;
	else
	if(re)				gb <=  1'b0;
 
////////////////////////////////////////////////////////////////////
//
// Registered Full & Empty Flags
//
 
// Guard Bit ...
always @(posedge clk )
	if(!rst)			gb2 <=  1'b0;
	else
	if(clr)				gb2 <=  1'b0;
	else
	if((wp_pl2 == rp) & we)		gb2 <=  1'b1;
	else
	if((wp != rp) & re)		gb2 <=  1'b0;
 
always @(posedge clk )
	if(!rst)				full_r <=  1'b0;
	else
	if(clr)					full_r <=  1'b0;
	else
	if(we & ((wp_pl1 == rp) & gb2) & !re)	full_r <=  1'b1;
	else
	if(re & ((wp_pl1 != rp) | !gb2) & !we)	full_r <=  1'b0;
 
always @(posedge clk )
	if(!rst)				empty_r <=  1'b1;
	else
	if(clr)					empty_r <=  1'b1;
	else
	if(we & ((wp != rp_pl1) | gb2) & !re)	empty_r <=  1'b0;
	else
	if(re & ((wp == rp_pl1) & !gb2) & !we)	empty_r <=  1'b1;
 
////////////////////////////////////////////////////////////////////
//
// Combinatorial Full_n & Empty_n Flags
//
 
assign empty_n = cnt < `n;
assign full_n  = !(cnt < (`max_size-`n+1));
assign level = {{cnt[`awa]}, {cnt[`awa]}} | cnt[`awa-1:`awa-2];
 
// N entries status
always @(posedge clk )
	if(!rst)	cnt <=  {4'b0000};
	else
	if(clr)		cnt <=  {4'b0000};
	else
	if( re & !we)	cnt <=  cnt + { 5'b11111};
	else
	if(!re &  we)	cnt <=  cnt + { {4'b0000}, 1'b1};
 
////////////////////////////////////////////////////////////////////
//
// Registered Full_n & Empty_n Flags
//
 
always @(posedge clk )
	if(!rst)				empty_n_r <=  1'b1;
	else
	if(clr)					empty_n_r <=  1'b1;
	else
	if(we & (cnt >= (`n-1) ) & !re)		empty_n_r <=  1'b0;
	else
	if(re & (cnt <= `n ) & !we)		empty_n_r <=  1'b1;
 
always @(posedge clk )
	if(!rst)				full_n_r <=  1'b0;
	else
	if(clr)					full_n_r <=  1'b0;
	else
	if(we & (cnt >= (`max_size-`n) ) & !re)	full_n_r <=  1'b1;
	else
	if(re & (cnt <= (`max_size-`n+1)) & !we)	full_n_r <=  1'b0;

endmodule
 

 
 
  
module arSRLFIFO_d (CLK, RST_N, D_IN,ENQ,DEQ,CLR,D_OUT,EMPTY_N,FULL_N);

input CLK;
input RST_N;
input [127:0] D_IN;
input ENQ;
input DEQ;
input CLR;
output [127:0] D_OUT;
output EMPTY_N;
output FULL_N;



wire fulln;
wire emptyn;

wire always_one;
wire always_zero;

assign always_one = 1'b1;
assign always_zero = 1'b0;

generic_fifo_sc_d fifo_1
(.clk(CLK),
 .rst(RST_N),
 .clr (CLR),
 .din (D_IN),
 .we (ENQ),
 .dout (D_OUT),
 .re (DEQ),
 .full_r (FULL_N),
 .empty_r(EMPTY_N),
 .full_n_r (fulln),
 .empty_n_r (emptyn)
 );
 







endmodule








/////////////////////////////////////////////////////////////////////
////                                                             ////
////  Universal FIFO Single Clock                                ////
////                                                             ////
////                                                             ////
////  Author: Rudolf Usselmann                                   ////
////          rudi@asics.ws                                      ////
////                                                             ////
////                                                             ////
////  D/L from: http://www.opencores.org/cores/generic_fifos/    ////
////                                                             ////
/////////////////////////////////////////////////////////////////////
////                                                             ////
//// Copyright (C) 2000-2002 Rudolf Usselmann                    ////
////                         www.asics.ws                        ////
////                         rudi@asics.ws                       ////
////                                                             ////
//// This source file may be used and distributed without        ////
//// restriction provided that this copyright statement is not   ////
//// removed from the file and that any derivative work contains ////
//// the original copyright notice and the associated disclaimer.////
////                                                             ////
////     THIS SOFTWARE IS PROVIDED ``AS IS'' AND WITHOUT ANY     ////
//// EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED   ////
//// TO, THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS   ////
//// FOR A PARTICULAR PURPOSE. IN NO EVENT SHALL THE AUTHOR      ////
//// OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT, INDIRECT,         ////
//// INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES    ////
//// (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE   ////
//// GOODS OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR        ////
//// BUSINESS INTERRUPTION) HOWEVER CAUSED AND ON ANY THEORY OF  ////
//// LIABILITY, WHETHER IN  CONTRACT, STRICT LIABILITY, OR TORT  ////
//// (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT  ////
//// OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED OF THE         ////
//// POSSIBILITY OF SUCH DAMAGE.                                 ////
////                                                             ////
/////////////////////////////////////////////////////////////////////
 
//  CVS Log
//
//  __Id: generic_fifo_sc_a.v,v 1.1.1.1 2002-09-25 05:42:06 rudi Exp __
//
//  __Date: 2002-09-25 05:42:06 __
//  __Revision: 1.1.1.1 __
//  __Author: rudi __
//  __Locker:  __
//  __State: Exp __
//
// Change History:
//               __Log: not supported by cvs2svn __
//
//
//
//
//
//
//
//
//
//
 
 
/*
 
Description
===========
 
I/Os
----
rst	low active, either sync. or async. master reset (see below how to select)
clr	synchronous clear (just like reset but always synchronous), high active
re	read enable, synchronous, high active
we	read enable, synchronous, high active
din	Data Input
dout	Data Output
 
full	Indicates the FIFO is full (combinatorial output)
full_r	same as above, but registered output (see note below)
empty	Indicates the FIFO is empty
empty_r	same as above, but registered output (see note below)
 
full_n		Indicates if the FIFO has space for N entries (combinatorial output)
full_n_r	same as above, but registered output (see note below)
empty_n		Indicates the FIFO has at least N entries (combinatorial output)
empty_n_r	same as above, but registered output (see note below)
 
level		indicates the FIFO level:
		2'b00	0-25%	 full
		2'b01	25-50%	 full
		2'b10	50-75%	 full
		2'b11	%75-100% full
 
combinatorial vs. registered status outputs
-------------------------------------------
Both the combinatorial and registered status outputs have exactly the same
synchronous timing. Meaning they are being asserted immediately at the clock
edge after the last read or write. The combinatorial outputs however, pass
through several levels of logic before they are output. The registered status
outputs are direct outputs of a flip-flop. The reason both are provided, is
that the registered outputs require quite a bit of additional logic inside
the FIFO. If you can meet timing of your device with the combinatorial
outputs, use them ! The FIFO will be smaller. If the status signals are
in the critical pass, use the registered outputs, they have a much smaller
output delay (actually only Tcq).
 
Parameters
----------
The FIFO takes 3 parameters:
dw	Data bus width
aw	Address bus width (Determines the FIFO size by evaluating 2^aw)
n	N is a second status threshold constant for full_n and empty_n
	If you have no need for the second status threshold, do not
	connect the outputs and the logic should be removed by your
	synthesis tool.
 
Synthesis Results
-----------------
In a Spartan 2e a 8 bit wide, 8 entries deep FIFO, takes 85 LUTs and runs
at about 116 MHz (IO insertion disabled). The registered status outputs
are valid after 2.1NS, the combinatorial once take out to 6.5 NS to be
available.
 
 
Misc
----
This design assumes you will do appropriate status checking externally.
 
IMPORTANT ! writing while the FIFO is full or reading while the FIFO is
empty will place the FIFO in an undefined state.
 
*/
 
 
// Selecting Sync. or Async Reset
// ------------------------------
// Uncomment one of the two lines below. The first line for
// synchronous reset, the second for asynchronous reset
 
//`define SC_FIFO_ASYNC_RESET				// Uncomment for Syncr. reset
//`define SC_FIFO_ASYNC_RESET	or negedge rst		// Uncomment for Async. reset

/*
parameter dw=8;
parameter aw=8;
parameter n=32;
parameter max_size = 1<<aw;
 */
 
 `define dwd 128 

module generic_fifo_sc_d(clk, rst, clr, din, we, dout, re,
			 full_r, empty_r,
			 full_n_r, empty_n_r);
 /*
parameter dw=8;
parameter aw=8;
parameter n=32;
parameter max_size = 1<<aw;
 */
input			clk, rst, clr;
input	[`dwd-1:0]	din;
input			we;
output	[`dwd-1:0]	dout;
input			re;
wire			full; output full_r;
wire			empty; output empty_r;
wire			full_n; output full_n_r;
wire			empty_n; output empty_n_r;
wire	[1:0]		level;
 
////////////////////////////////////////////////////////////////////
//
// Local Wires
//
 
reg	[`awa-1:0]	wp;
wire	[`awa-1:0]	wp_pl1;
wire	[`awa-1:0]	wp_pl2;
reg	[`awa-1:0]	rp;
wire	[`awa-1:0]	rp_pl1;
reg			full_r;
reg			empty_r;
reg			gb;
reg			gb2;
reg	[`awa:0]		cnt;
wire			full_n, empty_n;
reg			full_n_r, empty_n_r;
 
////////////////////////////////////////////////////////////////////
//
// Memory Block
//
 wire always_zero;
 assign always_zero = 1'b0;
 wire [`dwd-1:0] junk_out;
 
 wire [`dwd-1:0] junk_in;
 
 // manually assign
 assign junk_in = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
 
dual_port_ram   #( .ADDR_WIDTH(4), .DATA_WIDTH(128))  ram1(
	.clk(		clk		),
	.addr1(		rp		),
	.addr2(		wp		),
	.we1(		we		),
	.we2(		always_zero		),
	.out1(		dout		),
	.out2(		junk_out		),
	.data1(		din		),
	.data2 (	junk_in)
	);
 
////////////////////////////////////////////////////////////////////
//
// Misc Logic
//
 
always @(posedge clk )
	if(!rst)	wp <=  {4'b0000};
	else
	if(clr)		wp <=  {4'b0000};
	else
	if(we)		wp <=  wp_pl1;
 
assign wp_pl1 = wp + { {3'b000}, 1'b1};
assign wp_pl2 = wp + { {2'b00}, 2'b10};
 
always @(posedge clk )
	if(!rst)	rp <=  {4'b0000};
	else
	if(clr)		rp <=  {4'b0000};
	else
	if(re)		rp <=  rp_pl1;
 
assign rp_pl1 = rp + { {3'b000}, 1'b1};
 
////////////////////////////////////////////////////////////////////
//
// Combinatorial Full & Empty Flags
//
 
assign empty = ((wp == rp) & !gb);
assign full  = ((wp == rp) &  gb);
 
// Guard Bit ...
always @(posedge clk )
	if(!rst)			gb <=  1'b0;
	else
	if(clr)				gb <=  1'b0;
	else
	if((wp_pl1 == rp) & we)		gb <=  1'b1;
	else
	if(re)				gb <=  1'b0;
 
////////////////////////////////////////////////////////////////////
//
// Registered Full & Empty Flags
//
 
// Guard Bit ...
always @(posedge clk )
	if(!rst)			gb2 <=  1'b0;
	else
	if(clr)				gb2 <=  1'b0;
	else
	if((wp_pl2 == rp) & we)		gb2 <=  1'b1;
	else
	if((wp != rp) & re)		gb2 <=  1'b0;
 
always @(posedge clk )
	if(!rst)				full_r <=  1'b0;
	else
	if(clr)					full_r <=  1'b0;
	else
	if(we & ((wp_pl1 == rp) & gb2) & !re)	full_r <=  1'b1;
	else
	if(re & ((wp_pl1 != rp) | !gb2) & !we)	full_r <=  1'b0;
 
always @(posedge clk )
	if(!rst)				empty_r <=  1'b1;
	else
	if(clr)					empty_r <=  1'b1;
	else
	if(we & ((wp != rp_pl1) | gb2) & !re)	empty_r <=  1'b0;
	else
	if(re & ((wp == rp_pl1) & !gb2) & !we)	empty_r <=  1'b1;
 
////////////////////////////////////////////////////////////////////
//
// Combinatorial Full_n & Empty_n Flags
//
 
assign empty_n = cnt < `n;
assign full_n  = !(cnt < (`max_size-`n+1));
assign level = {{cnt[`awa]}, {cnt[`awa]}} | cnt[`awa-1:`awa-2];
 
// N entries status
always @(posedge clk )
	if(!rst)	cnt <=  {4'b0000};
	else
	if(clr)		cnt <=  {4'b0000};
	else
	if( re & !we)	cnt <=  cnt + { 5'b11111};
	else
	if(!re &  we)	cnt <=  cnt + { {4'b0000}, 1'b1};
 
////////////////////////////////////////////////////////////////////
//
// Registered Full_n & Empty_n Flags
//
 
always @(posedge clk )
	if(!rst)				empty_n_r <=  1'b1;
	else
	if(clr)					empty_n_r <=  1'b1;
	else
	if(we & (cnt >= (`n-1) ) & !re)		empty_n_r <=  1'b0;
	else
	if(re & (cnt <= `n ) & !we)		empty_n_r <=  1'b1;
 
always @(posedge clk )
	if(!rst)				full_n_r <=  1'b0;
	else
	if(clr)					full_n_r <=  1'b0;
	else
	if(we & (cnt >= (`max_size-`n) ) & !re)	full_n_r <=  1'b1;
	else
	if(re & (cnt <= (`max_size-`n+1)) & !we)	full_n_r <=  1'b0;

endmodule
 

 
 
module SizedFIFO_a (CLK, D_IN,ENQ,DEQ,CLR,D_OUT,FULL_N,EMPTY_N);


input CLK;
input [59:0] D_IN;
input ENQ;
input DEQ;
input	CLR;
output [59:0]	D_OUT;
output	FULL_N;
output	EMPTY_N;
		



wire fulln;
wire emptyn;

wire always_one;
wire always_zero;

assign always_one = 1'b1;
assign always_zero = 1'b0;

generic_fifo_sc_f fifo_1
(.clk(CLK),
 .rst(always_one),
 .clr (CLR),
 .din (D_IN),
 .we (ENQ),
 .dout (D_OUT),
 .re (DEQ),
 .full_r (FULL_N),
 .empty_r(EMPTY_N),
 .full_n_r (fulln),
 .empty_n_r (emptyn)
 );
 







endmodule








/////////////////////////////////////////////////////////////////////
////                                                             ////
////  Universal FIFO Single Clock                                ////
////                                                             ////
////                                                             ////
////  Author: Rudolf Usselmann                                   ////
////          rudi@asics.ws                                      ////
////                                                             ////
////                                                             ////
////  D/L from: http://www.opencores.org/cores/generic_fifos/    ////
////                                                             ////
/////////////////////////////////////////////////////////////////////
////                                                             ////
//// Copyright (C) 2000-2002 Rudolf Usselmann                    ////
////                         www.asics.ws                        ////
////                         rudi@asics.ws                       ////
////                                                             ////
//// This source file may be used and distributed without        ////
//// restriction provided that this copyright statement is not   ////
//// removed from the file and that any derivative work contains ////
//// the original copyright notice and the associated disclaimer.////
////                                                             ////
////     THIS SOFTWARE IS PROVIDED ``AS IS'' AND WITHOUT ANY     ////
//// EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED   ////
//// TO, THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS   ////
//// FOR A PARTICULAR PURPOSE. IN NO EVENT SHALL THE AUTHOR      ////
//// OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT, INDIRECT,         ////
//// INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES    ////
//// (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE   ////
//// GOODS OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR        ////
//// BUSINESS INTERRUPTION) HOWEVER CAUSED AND ON ANY THEORY OF  ////
//// LIABILITY, WHETHER IN  CONTRACT, STRICT LIABILITY, OR TORT  ////
//// (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT  ////
//// OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED OF THE         ////
//// POSSIBILITY OF SUCH DAMAGE.                                 ////
////                                                             ////
/////////////////////////////////////////////////////////////////////
 
//  CVS Log
//
//  __Id: generic_fifo_sc_a.v,v 1.1.1.1 2002-09-25 05:42:06 rudi Exp __
//
//  __Date: 2002-09-25 05:42:06 __
//  __Revision: 1.1.1.1 __
//  __Author: rudi __
//  __Locker:  __
//  __State: Exp __
//
// Change History:
//               __Log: not supported by cvs2svn __
//
//
//
//
//
//
//
//
//
//
 
 
/*
 
Description
===========
 
I/Os
----
rst	low active, either sync. or async. master reset (see below how to select)
clr	synchronous clear (just like reset but always synchronous), high active
re	read enable, synchronous, high active
we	read enable, synchronous, high active
din	Data Input
dout	Data Output
 
full	Indicates the FIFO is full (combinatorial output)
full_r	same as above, but registered output (see note below)
empty	Indicates the FIFO is empty
empty_r	same as above, but registered output (see note below)
 
full_n		Indicates if the FIFO has space for N entries (combinatorial output)
full_n_r	same as above, but registered output (see note below)
empty_n		Indicates the FIFO has at least N entries (combinatorial output)
empty_n_r	same as above, but registered output (see note below)
 
level		indicates the FIFO level:
		2'b00	0-25%	 full
		2'b01	25-50%	 full
		2'b10	50-75%	 full
		2'b11	%75-100% full
 
combinatorial vs. registered status outputs
-------------------------------------------
Both the combinatorial and registered status outputs have exactly the same
synchronous timing. Meaning they are being asserted immediately at the clock
edge after the last read or write. The combinatorial outputs however, pass
through several levels of logic before they are output. The registered status
outputs are direct outputs of a flip-flop. The reason both are provided, is
that the registered outputs require quite a bit of additional logic inside
the FIFO. If you can meet timing of your device with the combinatorial
outputs, use them ! The FIFO will be smaller. If the status signals are
in the critical pass, use the registered outputs, they have a much smaller
output delay (actually only Tcq).
 
Parameters
----------
The FIFO takes 3 parameters:
dw	Data bus width
aw	Address bus width (Determines the FIFO size by evaluating 2^aw)
n	N is a second status threshold constant for full_n and empty_n
	If you have no need for the second status threshold, do not
	connect the outputs and the logic should be removed by your
	synthesis tool.
 
Synthesis Results
-----------------
In a Spartan 2e a 8 bit wide, 8 entries deep FIFO, takes 85 LUTs and runs
at about 116 MHz (IO insertion disabled). The registered status outputs
are valid after 2.1NS, the combinatorial once take out to 6.5 NS to be
available.
 
 
Misc
----
This design assumes you will do appropriate status checking externally.
 
IMPORTANT ! writing while the FIFO is full or reading while the FIFO is
empty will place the FIFO in an undefined state.
 
*/
 
 
// Selecting Sync. or Async Reset
// ------------------------------
// Uncomment one of the two lines below. The first line for
// synchronous reset, the second for asynchronous reset
 
//`define SC_FIFO_ASYNC_RESET				// Uncomment for Syncr. reset
//`define SC_FIFO_ASYNC_RESET	or negedge rst		// Uncomment for Async. reset

/*
parameter dw=8;
parameter aw=8;
parameter n=32;
parameter max_size = 1<<aw;
 */
 
 `define dwc  60
`define awc 3

module generic_fifo_sc_f(clk, rst, clr, din, we, dout, re,
			 full_r, empty_r,
			 full_n_r, empty_n_r);
 /*
parameter dw=8;
parameter aw=8;
parameter n=32;
parameter max_size = 1<<aw;
 */
input			clk, rst, clr;
input	[`dwc-1:0]	din;
input			we;
output	[`dwc-1:0]	dout;
input			re;
wire			full; output full_r;
wire			empty; output empty_r;
wire			full_n; output full_n_r;
wire			empty_n; output empty_n_r;
wire	[1:0]		level;
 
////////////////////////////////////////////////////////////////////
//
// Local Wires
//
 
reg	[`awc-1:0]	wp;
wire	[`awc-1:0]	wp_pl1;
wire	[`awc-1:0]	wp_pl2;
reg	[`awc-1:0]	rp;
wire	[`awc-1:0]	rp_pl1;
reg			full_r;
reg			empty_r;
reg			gb;
reg			gb2;
reg	[`awc:0]		cnt;
wire			full_n, empty_n;
reg			full_n_r, empty_n_r;
 
////////////////////////////////////////////////////////////////////
//
// Memory Block
//
 wire always_zero;
 assign always_zero = 1'b0;
 wire [`dwc-1:0] junk_out;
 
 wire [`dwc-1:0] junk_in;
 
 // manually assign
 assign junk_in = 60'b000000000000000000000000000000000000000000000000000000000000;
 
dual_port_ram  #( .ADDR_WIDTH(4), .DATA_WIDTH(60))   ram1(
	.clk(		clk		),
	.addr1(		rp		),
	.addr2(		wp		),
	.we1(		we		),
	.we2(		always_zero		),
	.out1(		dout		),
	.out2(		junk_out		),
	.data1(		din		),
	.data2 (	junk_in)
	);
 
////////////////////////////////////////////////////////////////////
//
// Misc Logic
//
 
always @(posedge clk )
	if(!rst)	wp <=  {3'b000};
	else
	if(clr)		wp <=  {3'b000};
	else
	if(we)		wp <=  wp_pl1;
 
assign wp_pl1 = wp + { {2'b00}, 1'b1};
assign wp_pl2 = wp +  { {1'b0}, 2'b10};
 
always @(posedge clk )
	if(!rst)	rp <=  {3'b000};
	else
	if(clr)		rp <=  {3'b000};
	else
	if(re)		rp <=  rp_pl1;
 
assign rp_pl1 = rp + { {2'b00}, 1'b1};
 
////////////////////////////////////////////////////////////////////
//
// Combinatorial Full & Empty Flags
//
 
assign empty = ((wp == rp) & !gb);
assign full  = ((wp == rp) &  gb);
 
// Guard Bit ...
always @(posedge clk )
	if(!rst)			gb <=  1'b0;
	else
	if(clr)				gb <=  1'b0;
	else
	if((wp_pl1 == rp) & we)		gb <=  1'b1;
	else
	if(re)				gb <=  1'b0;
 
////////////////////////////////////////////////////////////////////
//
// Registered Full & Empty Flags
//
 
// Guard Bit ...
always @(posedge clk )
	if(!rst)			gb2 <=  1'b0;
	else
	if(clr)				gb2 <=  1'b0;
	else
	if((wp_pl2 == rp) & we)		gb2 <=  1'b1;
	else
	if((wp != rp) & re)		gb2 <=  1'b0;
 
always @(posedge clk )
	if(!rst)				full_r <=  1'b0;
	else
	if(clr)					full_r <=  1'b0;
	else
	if(we & ((wp_pl1 == rp) & gb2) & !re)	full_r <=  1'b1;
	else
	if(re & ((wp_pl1 != rp) | !gb2) & !we)	full_r <=  1'b0;
 
always @(posedge clk )
	if(!rst)				empty_r <=  1'b1;
	else
	if(clr)					empty_r <=  1'b1;
	else
	if(we & ((wp != rp_pl1) | gb2) & !re)	empty_r <=  1'b0;
	else
	if(re & ((wp == rp_pl1) & !gb2) & !we)	empty_r <=  1'b1;
 
////////////////////////////////////////////////////////////////////
//
// Combinatorial Full_n & Empty_n Flags
//
 
assign empty_n = cnt < `n;
assign full_n  = !(cnt < (`max_size-`n+1));
assign level = {{cnt[`awc]}, {cnt[`awc]}} | cnt[`awc-1:`awc-2];
 
// N entries status
always @(posedge clk )
	if(!rst)	cnt <=  {4'b0000};
	else
	if(clr)		cnt <=  {4'b0000};
	else
	if( re & !we)	cnt <=  cnt + { 4'b1111};
	else
	if(!re &  we)	cnt <=  cnt + { {3'b000}, 1'b1};
 
////////////////////////////////////////////////////////////////////
//
// Registered Full_n & Empty_n Flags
//
 
always @(posedge clk )
	if(!rst)				empty_n_r <=  1'b1;
	else
	if(clr)					empty_n_r <=  1'b1;
	else
	if(we & (cnt >= (`n-1) ) & !re)		empty_n_r <=  1'b0;
	else
	if(re & (cnt <= `n ) & !we)		empty_n_r <=  1'b1;
 
always @(posedge clk )
	if(!rst)				full_n_r <=  1'b0;
	else
	if(clr)					full_n_r <=  1'b0;
	else
	if(we & (cnt >= (`max_size-`n) ) & !re)	full_n_r <=  1'b1;
	else
	if(re & (cnt <= (`max_size-`n+1)) & !we)	full_n_r <=  1'b0;

endmodule
 
module SizedFIFO_b (CLK, D_IN,ENQ,DEQ,CLR,D_OUT,FULL_N,EMPTY_N);


input CLK;
input [312:0] D_IN;
input ENQ;
input DEQ;
input	CLR;
output [312:0]	D_OUT;
output	FULL_N;
output	EMPTY_N;
		



wire fulln;
wire emptyn;

wire always_one;
wire always_zero;

assign always_one = 1'b1;
assign always_zero = 1'b0;

generic_fifo_sc_g fifo_1
(.clk(CLK),
 .rst(always_one),
 .clr (CLR),
 .din (D_IN),
 .we (ENQ),
 .dout (D_OUT),
 .re (DEQ),
 .full_r (FULL_N),
 .empty_r(EMPTY_N),
 .full_n_r (fulln),
 .empty_n_r (emptyn)
 );
 







endmodule








/////////////////////////////////////////////////////////////////////
////                                                             ////
////  Universal FIFO Single Clock                                ////
////                                                             ////
////                                                             ////
////  Author: Rudolf Usselmann                                   ////
////          rudi@asics.ws                                      ////
////                                                             ////
////                                                             ////
////  D/L from: http://www.opencores.org/cores/generic_fifos/    ////
////                                                             ////
/////////////////////////////////////////////////////////////////////
////                                                             ////
//// Copyright (C) 2000-2002 Rudolf Usselmann                    ////
////                         www.asics.ws                        ////
////                         rudi@asics.ws                       ////
////                                                             ////
//// This source file may be used and distributed without        ////
//// restriction provided that this copyright statement is not   ////
//// removed from the file and that any derivative work contains ////
//// the original copyright notice and the associated disclaimer.////
////                                                             ////
////     THIS SOFTWARE IS PROVIDED ``AS IS'' AND WITHOUT ANY     ////
//// EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED   ////
//// TO, THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS   ////
//// FOR A PARTICULAR PURPOSE. IN NO EVENT SHALL THE AUTHOR      ////
//// OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT, INDIRECT,         ////
//// INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES    ////
//// (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE   ////
//// GOODS OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR        ////
//// BUSINESS INTERRUPTION) HOWEVER CAUSED AND ON ANY THEORY OF  ////
//// LIABILITY, WHETHER IN  CONTRACT, STRICT LIABILITY, OR TORT  ////
//// (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT  ////
//// OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED OF THE         ////
//// POSSIBILITY OF SUCH DAMAGE.                                 ////
////                                                             ////
/////////////////////////////////////////////////////////////////////
 
//  CVS Log
//
//  __Id: generic_fifo_sc_a.v,v 1.1.1.1 2002-09-25 05:42:06 rudi Exp __
//
//  __Date: 2002-09-25 05:42:06 __
//  __Revision: 1.1.1.1 __
//  __Author: rudi __
//  __Locker:  __
//  __State: Exp __
//
// Change History:
//               __Log: not supported by cvs2svn __
//
//
//
//
//
//
//
//
//
//
 
 
/*
 
Description
===========
 
I/Os
----
rst	low active, either sync. or async. master reset (see below how to select)
clr	synchronous clear (just like reset but always synchronous), high active
re	read enable, synchronous, high active
we	read enable, synchronous, high active
din	Data Input
dout	Data Output
 
full	Indicates the FIFO is full (combinatorial output)
full_r	same as above, but registered output (see note below)
empty	Indicates the FIFO is empty
empty_r	same as above, but registered output (see note below)
 
full_n		Indicates if the FIFO has space for N entries (combinatorial output)
full_n_r	same as above, but registered output (see note below)
empty_n		Indicates the FIFO has at least N entries (combinatorial output)
empty_n_r	same as above, but registered output (see note below)
 
level		indicates the FIFO level:
		2'b00	0-25%	 full
		2'b01	25-50%	 full
		2'b10	50-75%	 full
		2'b11	%75-100% full
 
combinatorial vs. registered status outputs
-------------------------------------------
Both the combinatorial and registered status outputs have exactly the same
synchronous timing. Meaning they are being asserted immediately at the clock
edge after the last read or write. The combinatorial outputs however, pass
through several levels of logic before they are output. The registered status
outputs are direct outputs of a flip-flop. The reason both are provided, is
that the registered outputs require quite a bit of additional logic inside
the FIFO. If you can meet timing of your device with the combinatorial
outputs, use them ! The FIFO will be smaller. If the status signals are
in the critical pass, use the registered outputs, they have a much smaller
output delay (actually only Tcq).
 
Parameters
----------
The FIFO takes 3 parameters:
dw	Data bus width
aw	Address bus width (Determines the FIFO size by evaluating 2^aw)
n	N is a second status threshold constant for full_n and empty_n
	If you have no need for the second status threshold, do not
	connect the outputs and the logic should be removed by your
	synthesis tool.
 
Synthesis Results
-----------------
In a Spartan 2e a 8 bit wide, 8 entries deep FIFO, takes 85 LUTs and runs
at about 116 MHz (IO insertion disabled). The registered status outputs
are valid after 2.1NS, the combinatorial once take out to 6.5 NS to be
available.
 
 
Misc
----
This design assumes you will do appropriate status checking externally.
 
IMPORTANT ! writing while the FIFO is full or reading while the FIFO is
empty will place the FIFO in an undefined state.
 
*/
 
 
// Selecting Sync. or Async Reset
// ------------------------------
// Uncomment one of the two lines below. The first line for
// synchronous reset, the second for asynchronous reset
 
//`define SC_FIFO_ASYNC_RESET				// Uncomment for Syncr. reset
//`define SC_FIFO_ASYNC_RESET	or negedge rst		// Uncomment for Async. reset

/*
parameter dw=8;
parameter aw=8;
parameter n=32;
parameter max_size = 1<<aw;
 */
 
 `define dwf  313
`define awf 3

module generic_fifo_sc_g(clk, rst, clr, din, we, dout, re,
			 full_r, empty_r,
			 full_n_r, empty_n_r);
 /*
parameter dw=8;
parameter aw=8;
parameter n=32;
parameter max_size = 1<<aw;
 */
input			clk, rst, clr;
input	[`dwf-1:0]	din;
input			we;
output	[`dwf-1:0]	dout;
input			re;
wire			full; output full_r;
wire			empty; output empty_r;
wire			full_n; output full_n_r;
wire			empty_n; output empty_n_r;
wire	[1:0]		level;
 
////////////////////////////////////////////////////////////////////
//
// Local Wires
//
 
reg	[`awf-1:0]	wp;
wire	[`awf-1:0]	wp_pl1;
wire	[`awf-1:0]	wp_pl2;
reg	[`awf-1:0]	rp;
wire	[`awf-1:0]	rp_pl1;
reg			full_r;
reg			empty_r;
reg			gb;
reg			gb2;
reg	[`awf:0]		cnt;
wire			full_n, empty_n;
reg			full_n_r, empty_n_r;
 
////////////////////////////////////////////////////////////////////
//
// Memory Block
//
 wire always_zero;
 assign always_zero = 1'b0;
 wire [`dwf-1:0] junk_out;
 
 wire [`dwf-1:0] junk_in;
 
 // manually assign
 assign junk_in = 313'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
 
dual_port_ram   #( .ADDR_WIDTH(4), .DATA_WIDTH(313))  ram1(
	.clk(		clk		),
	.addr1(		rp		),
	.addr2(		wp		),
	.we1(		we		),
	.we2(		always_zero		),
	.out1(		dout		),
	.out2(		junk_out		),
	.data1(		din		),
	.data2 (	junk_in)
	);
 
////////////////////////////////////////////////////////////////////
//
// Misc Logic
//
 
always @(posedge clk )
	if(!rst)	wp <=  {3'b000};
	else
	if(clr)		wp <=  {3'b000};
	else
	if(we)		wp <=  wp_pl1;
 
assign wp_pl1 = wp + { {2'b00}, 1'b1};
assign wp_pl2 = wp +  { {1'b0}, 2'b10};
 
always @(posedge clk )
	if(!rst)	rp <=  {3'b000};
	else
	if(clr)		rp <=  {3'b000};
	else
	if(re)		rp <=  rp_pl1;
 
assign rp_pl1 = rp + { {2'b00}, 1'b1};
 
////////////////////////////////////////////////////////////////////
//
// Combinatorial Full & Empty Flags
//
 
assign empty = ((wp == rp) & !gb);
assign full  = ((wp == rp) &  gb);
 
// Guard Bit ...
always @(posedge clk )
	if(!rst)			gb <=  1'b0;
	else
	if(clr)				gb <=  1'b0;
	else
	if((wp_pl1 == rp) & we)		gb <=  1'b1;
	else
	if(re)				gb <=  1'b0;
 
////////////////////////////////////////////////////////////////////
//
// Registered Full & Empty Flags
//
 
// Guard Bit ...
always @(posedge clk )
	if(!rst)			gb2 <=  1'b0;
	else
	if(clr)				gb2 <=  1'b0;
	else
	if((wp_pl2 == rp) & we)		gb2 <=  1'b1;
	else
	if((wp != rp) & re)		gb2 <=  1'b0;
 
always @(posedge clk )
	if(!rst)				full_r <=  1'b0;
	else
	if(clr)					full_r <=  1'b0;
	else
	if(we & ((wp_pl1 == rp) & gb2) & !re)	full_r <=  1'b1;
	else
	if(re & ((wp_pl1 != rp) | !gb2) & !we)	full_r <=  1'b0;
 
always @(posedge clk )
	if(!rst)				empty_r <=  1'b1;
	else
	if(clr)					empty_r <=  1'b1;
	else
	if(we & ((wp != rp_pl1) | gb2) & !re)	empty_r <=  1'b0;
	else
	if(re & ((wp == rp_pl1) & !gb2) & !we)	empty_r <=  1'b1;
 
////////////////////////////////////////////////////////////////////
//
// Combinatorial Full_n & Empty_n Flags
//
 
assign empty_n = cnt < `n;
assign full_n  = !(cnt < (`max_size-`n+1));
assign level = {{cnt[`awf]}, {cnt[`awf]}} | cnt[`awf-1:`awf-2];
 
// N entries status
always @(posedge clk )
	if(!rst)	cnt <=  {3'b000};
	else
	if(clr)		cnt <=  {3'b000};
	else
	if( re & !we)	cnt <=  cnt + { 4'b1111};
	else
	if(!re &  we)	cnt <=  cnt + { {3'b000}, 1'b1};
 
////////////////////////////////////////////////////////////////////
//
// Registered Full_n & Empty_n Flags
//
 
always @(posedge clk )
	if(!rst)				empty_n_r <=  1'b1;
	else
	if(clr)					empty_n_r <=  1'b1;
	else
	if(we & (cnt >= (`n-1) ) & !re)		empty_n_r <=  1'b0;
	else
	if(re & (cnt <= `n ) & !we)		empty_n_r <=  1'b1;
 
always @(posedge clk )
	if(!rst)				full_n_r <=  1'b0;
	else
	if(clr)					full_n_r <=  1'b0;
	else
	if(we & (cnt >= (`max_size-`n) ) & !re)	full_n_r <=  1'b1;
	else
	if(re & (cnt <= (`max_size-`n+1)) & !we)	full_n_r <=  1'b0;

endmodule




module SizedFIFO_x (CLK, D_IN,ENQ,DEQ,CLR,D_OUT,FULL_N,EMPTY_N);


input CLK;
input [130:0] D_IN;
input ENQ;
input DEQ;
input	CLR;
output [130:0]	D_OUT;
output	FULL_N;
output	EMPTY_N;
		



wire fulln;
wire emptyn;

wire always_one;
wire always_zero;

assign always_one = 1'b1;
assign always_zero = 1'b0;

generic_fifo_sc_x fifo_1
(.clk(CLK),
 .rst(always_one),
 .clr (CLR),
 .din (D_IN),
 .we (ENQ),
 .dout (D_OUT),
 .re (DEQ),
 .full_r (FULL_N),
 .empty_r(EMPTY_N),
 .full_n_r (fulln),
 .empty_n_r (emptyn)
 );
 







endmodule








/////////////////////////////////////////////////////////////////////
////                                                             ////
////  Universal FIFO Single Clock                                ////
////                                                             ////
////                                                             ////
////  Author: Rudolf Usselmann                                   ////
////          rudi@asics.ws                                      ////
////                                                             ////
////                                                             ////
////  D/L from: http://www.opencores.org/cores/generic_fifos/    ////
////                                                             ////
/////////////////////////////////////////////////////////////////////
////                                                             ////
//// Copyright (C) 2000-2002 Rudolf Usselmann                    ////
////                         www.asics.ws                        ////
////                         rudi@asics.ws                       ////
////                                                             ////
//// This source file may be used and distributed without        ////
//// restriction provided that this copyright statement is not   ////
//// removed from the file and that any derivative work contains ////
//// the original copyright notice and the associated disclaimer.////
////                                                             ////
////     THIS SOFTWARE IS PROVIDED ``AS IS'' AND WITHOUT ANY     ////
//// EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED   ////
//// TO, THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS   ////
//// FOR A PARTICULAR PURPOSE. IN NO EVENT SHALL THE AUTHOR      ////
//// OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT, INDIRECT,         ////
//// INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES    ////
//// (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE   ////
//// GOODS OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR        ////
//// BUSINESS INTERRUPTION) HOWEVER CAUSED AND ON ANY THEORY OF  ////
//// LIABILITY, WHETHER IN  CONTRACT, STRICT LIABILITY, OR TORT  ////
//// (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT  ////
//// OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED OF THE         ////
//// POSSIBILITY OF SUCH DAMAGE.                                 ////
////                                                             ////
/////////////////////////////////////////////////////////////////////
 
//  CVS Log
//
//  __Id: generic_fifo_sc_a.v,v 1.1.1.1 2002-09-25 05:42:06 rudi Exp __
//
//  __Date: 2002-09-25 05:42:06 __
//  __Revision: 1.1.1.1 __
//  __Author: rudi __
//  __Locker:  __
//  __State: Exp __
//
// Change History:
//               __Log: not supported by cvs2svn __
//
//
//
//
//
//
//
//
//
//
 
 
/*
 
Description
===========
 
I/Os
----
rst	low active, either sync. or async. master reset (see below how to select)
clr	synchronous clear (just like reset but always synchronous), high active
re	read enable, synchronous, high active
we	read enable, synchronous, high active
din	Data Input
dout	Data Output
 
full	Indicates the FIFO is full (combinatorial output)
full_r	same as above, but registered output (see note below)
empty	Indicates the FIFO is empty
empty_r	same as above, but registered output (see note below)
 
full_n		Indicates if the FIFO has space for N entries (combinatorial output)
full_n_r	same as above, but registered output (see note below)
empty_n		Indicates the FIFO has at least N entries (combinatorial output)
empty_n_r	same as above, but registered output (see note below)
 
level		indicates the FIFO level:
		2'b00	0-25%	 full
		2'b01	25-50%	 full
		2'b10	50-75%	 full
		2'b11	%75-100% full
 
combinatorial vs. registered status outputs
-------------------------------------------
Both the combinatorial and registered status outputs have exactly the same
synchronous timing. Meaning they are being asserted immediately at the clock
edge after the last read or write. The combinatorial outputs however, pass
through several levels of logic before they are output. The registered status
outputs are direct outputs of a flip-flop. The reason both are provided, is
that the registered outputs require quite a bit of additional logic inside
the FIFO. If you can meet timing of your device with the combinatorial
outputs, use them ! The FIFO will be smaller. If the status signals are
in the critical pass, use the registered outputs, they have a much smaller
output delay (actually only Tcq).
 
Parameters
----------
The FIFO takes 3 parameters:
dw	Data bus width
aw	Address bus width (Determines the FIFO size by evaluating 2^aw)
n	N is a second status threshold constant for full_n and empty_n
	If you have no need for the second status threshold, do not
	connect the outputs and the logic should be removed by your
	synthesis tool.
 
Synthesis Results
-----------------
In a Spartan 2e a 8 bit wide, 8 entries deep FIFO, takes 85 LUTs and runs
at about 116 MHz (IO insertion disabled). The registered status outputs
are valid after 2.1NS, the combinatorial once take out to 6.5 NS to be
available.
 
 
Misc
----
This design assumes you will do appropriate status checking externally.
 
IMPORTANT ! writing while the FIFO is full or reading while the FIFO is
empty will place the FIFO in an undefined state.
 
*/
 
 
// Selecting Sync. or Async Reset
// ------------------------------
// Uncomment one of the two lines below. The first line for
// synchronous reset, the second for asynchronous reset
 
//`define SC_FIFO_ASYNC_RESET				// Uncomment for Syncr. reset
//`define SC_FIFO_ASYNC_RESET	or negedge rst		// Uncomment for Async. reset

/*
parameter dw=8;
parameter aw=8;
parameter n=32;
parameter max_size = 1<<aw;
 */
 
 `define dwx  131
`define awx 2

module generic_fifo_sc_x(clk, rst, clr, din, we, dout, re,
			 full_r, empty_r,
			 full_n_r, empty_n_r);
 /*
parameter dw=8;
parameter aw=8;
parameter n=32;
parameter max_size = 1<<aw;
 */
input			clk, rst, clr;
input	[`dwx-1:0]	din;
input			we;
output	[`dwx-1:0]	dout;
input			re;
wire			full; output full_r;
wire			empty; output empty_r;
wire			full_n; output full_n_r;
wire			empty_n; output empty_n_r;
wire	[1:0]		level;
 
////////////////////////////////////////////////////////////////////
//
// Local Wires
//
 
reg	[`awx-1:0]	wp;
wire	[`awx-1:0]	wp_pl1;
wire	[`awx-1:0]	wp_pl2;
reg	[`awx-1:0]	rp;
wire	[`awx-1:0]	rp_pl1;
reg			full_r;
reg			empty_r;
reg			gb;
reg			gb2;
reg	[`awx:0]		cnt;
wire			full_n, empty_n;
reg			full_n_r, empty_n_r;
 
////////////////////////////////////////////////////////////////////
//
// Memory Block
//
 wire always_zero;
 assign always_zero = 1'b0;
 wire [`dwx-1:0] junk_out;
 
 wire [`dwx-1:0] junk_in;
 
 // manually assign
 assign junk_in = 131'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
 
dual_port_ram  #( .ADDR_WIDTH(4), .DATA_WIDTH(131))   ram1(
	.clk(		clk		),
	.addr1(		rp		),
	.addr2(		wp		),
	.we1(		we		),
	.we2(		always_zero		),
	.out1(		dout		),
	.out2(		junk_out		),
	.data1(		din		),
	.data2 (	junk_in)
	);
 
////////////////////////////////////////////////////////////////////
//
// Misc Logic
//
 
always @(posedge clk )
	if(!rst)	wp <=  {2'b00};
	else
	if(clr)		wp <=  {2'b00};
	else
	if(we)		wp <=  wp_pl1;
 
assign wp_pl1 = wp + { {1'b0}, 1'b1};
assign wp_pl2 = wp +  {  2'b10};
 
always @(posedge clk )
	if(!rst)	rp <=  {2'b00};
	else
	if(clr)		rp <=  {2'b00};
	else
	if(re)		rp <=  rp_pl1;
 
assign rp_pl1 = rp + { {1'b0}, 1'b1};
 
////////////////////////////////////////////////////////////////////
//
// Combinatorial Full & Empty Flags
//
 
assign empty = ((wp == rp) & !gb);
assign full  = ((wp == rp) &  gb);
 
// Guard Bit ...
always @(posedge clk )
	if(!rst)			gb <=  1'b0;
	else
	if(clr)				gb <=  1'b0;
	else
	if((wp_pl1 == rp) & we)		gb <=  1'b1;
	else
	if(re)				gb <=  1'b0;
 
////////////////////////////////////////////////////////////////////
//
// Registered Full & Empty Flags
//
 
// Guard Bit ...
always @(posedge clk )
	if(!rst)			gb2 <=  1'b0;
	else
	if(clr)				gb2 <=  1'b0;
	else
	if((wp_pl2 == rp) & we)		gb2 <=  1'b1;
	else
	if((wp != rp) & re)		gb2 <=  1'b0;
 
always @(posedge clk )
	if(!rst)				full_r <=  1'b0;
	else
	if(clr)					full_r <=  1'b0;
	else
	if(we & ((wp_pl1 == rp) & gb2) & !re)	full_r <=  1'b1;
	else
	if(re & ((wp_pl1 != rp) | !gb2) & !we)	full_r <=  1'b0;
 
always @(posedge clk )
	if(!rst)				empty_r <=  1'b1;
	else
	if(clr)					empty_r <=  1'b1;
	else
	if(we & ((wp != rp_pl1) | gb2) & !re)	empty_r <=  1'b0;
	else
	if(re & ((wp == rp_pl1) & !gb2) & !we)	empty_r <=  1'b1;
 
////////////////////////////////////////////////////////////////////
//
// Combinatorial Full_n & Empty_n Flags
//
 
assign empty_n = cnt < `n;
assign full_n  = !(cnt < (`max_size-`n+1));
assign level = {{cnt[`awx]}, {cnt[`awx]}} | cnt[`awx-1:`awx-2];
 
// N entries status
always @(posedge clk )
	if(!rst)	cnt <=  {3'b000};
	else
	if(clr)		cnt <=  {3'b000};
	else
	if( re & !we)	cnt <=  cnt + { 3'b1111};
	else
	if(!re &  we)	cnt <=  cnt + { {2'b00}, 1'b1};
 
////////////////////////////////////////////////////////////////////
//
// Registered Full_n & Empty_n Flags
//
 
always @(posedge clk )
	if(!rst)				empty_n_r <=  1'b1;
	else
	if(clr)					empty_n_r <=  1'b1;
	else
	if(we & (cnt >= (`n-1) ) & !re)		empty_n_r <=  1'b0;
	else
	if(re & (cnt <= `n ) & !we)		empty_n_r <=  1'b1;
 
always @(posedge clk )
	if(!rst)				full_n_r <=  1'b0;
	else
	if(clr)					full_n_r <=  1'b0;
	else
	if(we & (cnt >= (`max_size-`n) ) & !re)	full_n_r <=  1'b1;
	else
	if(re & (cnt <= (`max_size-`n+1)) & !we)	full_n_r <=  1'b0;

endmodule
